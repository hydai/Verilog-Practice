
module SingleCycleProcessor_DW_cmp_0 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, 
        EQ_NE );
  input [31:0] A;
  input [31:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325;

  OAI32XL U157 ( .A0(n262), .A1(A[2]), .A2(n314), .B0(A[3]), .B1(n261), .Y(
        n312) );
  OAI32XL U158 ( .A0(n252), .A1(A[20]), .A2(n275), .B0(A[21]), .B1(n251), .Y(
        n273) );
  NOR2BXL U159 ( .AN(A[21]), .B(B[21]), .Y(n275) );
  INVXL U160 ( .A(A[1]), .Y(n243) );
  AOI21XL U161 ( .A0(A[2]), .A1(n262), .B0(n314), .Y(n313) );
  AOI2BB1XL U162 ( .A0N(n243), .A1N(B[1]), .B0(A[0]), .Y(n311) );
  OAI211XL U163 ( .A0(B[12]), .A1(n235), .B0(n320), .C0(n318), .Y(n300) );
  AOI32XL U164 ( .A0(B[12]), .A1(n235), .A2(n320), .B0(n234), .B1(B[13]), .Y(
        n319) );
  NOR2BXL U165 ( .AN(A[7]), .B(B[7]), .Y(n310) );
  OR2XL U166 ( .A(B[11]), .B(n236), .Y(n324) );
  OR2XL U167 ( .A(B[9]), .B(n238), .Y(n302) );
  OAI32XL U168 ( .A0(n260), .A1(A[6]), .A2(n310), .B0(A[7]), .B1(n259), .Y(
        n309) );
  AOI32XL U169 ( .A0(B[8]), .A1(n239), .A2(n302), .B0(n238), .B1(B[9]), .Y(
        n323) );
  AOI32XL U170 ( .A0(B[10]), .A1(n237), .A2(n324), .B0(n236), .B1(B[11]), .Y(
        n322) );
  INVXL U171 ( .A(B[2]), .Y(n262) );
  INVXL U172 ( .A(B[6]), .Y(n260) );
  INVXL U173 ( .A(B[3]), .Y(n261) );
  INVXL U174 ( .A(B[7]), .Y(n259) );
  CLKINVX1 U175 ( .A(n282), .Y(n231) );
  CLKINVX1 U176 ( .A(n274), .Y(n232) );
  INVXL U177 ( .A(A[28]), .Y(n230) );
  INVXL U178 ( .A(A[29]), .Y(n229) );
  CLKINVX1 U179 ( .A(A[12]), .Y(n235) );
  CLKINVX1 U180 ( .A(A[4]), .Y(n242) );
  CLKINVX1 U181 ( .A(A[10]), .Y(n237) );
  CLKINVX1 U182 ( .A(A[8]), .Y(n239) );
  CLKINVX1 U183 ( .A(A[13]), .Y(n234) );
  CLKINVX1 U184 ( .A(A[11]), .Y(n236) );
  CLKINVX1 U185 ( .A(A[9]), .Y(n238) );
  CLKINVX1 U186 ( .A(A[5]), .Y(n241) );
  CLKINVX1 U187 ( .A(B[19]), .Y(n253) );
  CLKINVX1 U188 ( .A(B[21]), .Y(n251) );
  CLKINVX1 U189 ( .A(n288), .Y(n228) );
  CLKINVX1 U190 ( .A(A[31]), .Y(n227) );
  CLKINVX1 U191 ( .A(n319), .Y(n233) );
  CLKINVX1 U192 ( .A(B[15]), .Y(n257) );
  CLKINVX1 U193 ( .A(B[27]), .Y(n245) );
  CLKINVX1 U194 ( .A(B[25]), .Y(n247) );
  CLKINVX1 U195 ( .A(n309), .Y(n240) );
  CLKINVX1 U196 ( .A(B[14]), .Y(n258) );
  CLKINVX1 U197 ( .A(B[20]), .Y(n252) );
  CLKINVX1 U198 ( .A(B[24]), .Y(n248) );
  CLKINVX1 U199 ( .A(B[22]), .Y(n250) );
  CLKINVX1 U200 ( .A(B[18]), .Y(n254) );
  CLKINVX1 U201 ( .A(B[30]), .Y(n244) );
  CLKINVX1 U202 ( .A(B[26]), .Y(n246) );
  CLKINVX1 U203 ( .A(B[17]), .Y(n255) );
  CLKINVX1 U204 ( .A(B[23]), .Y(n249) );
  CLKINVX1 U205 ( .A(B[16]), .Y(n256) );
  OAI31XL U206 ( .A0(n263), .A1(n264), .A2(n265), .B0(n266), .Y(GE_LT_GT_LE)
         );
  OAI22XL U207 ( .A0(n267), .A1(n268), .B0(n269), .B1(n267), .Y(n266) );
  OAI21XL U208 ( .A0(n231), .A1(n270), .B0(n271), .Y(n268) );
  OAI22XL U209 ( .A0(n272), .A1(n273), .B0(n274), .B1(n272), .Y(n271) );
  OAI32X1 U210 ( .A0(n250), .A1(A[22]), .A2(n276), .B0(A[23]), .B1(n249), .Y(
        n272) );
  OAI22XL U211 ( .A0(n277), .A1(n278), .B0(n279), .B1(n277), .Y(n270) );
  OAI32X1 U212 ( .A0(n256), .A1(A[16]), .A2(n280), .B0(A[17]), .B1(n255), .Y(
        n278) );
  OAI32X1 U213 ( .A0(n254), .A1(A[18]), .A2(n281), .B0(A[19]), .B1(n253), .Y(
        n277) );
  OAI21XL U214 ( .A0(n283), .A1(n284), .B0(n285), .Y(n267) );
  OAI22XL U215 ( .A0(n286), .A1(n228), .B0(n287), .B1(n286), .Y(n285) );
  AOI32X1 U216 ( .A0(B[28]), .A1(n230), .A2(n289), .B0(n229), .B1(B[29]), .Y(
        n288) );
  OAI32X1 U217 ( .A0(n244), .A1(A[30]), .A2(n290), .B0(B[31]), .B1(n227), .Y(
        n286) );
  OAI22XL U218 ( .A0(n291), .A1(n292), .B0(n293), .B1(n291), .Y(n284) );
  OAI32X1 U219 ( .A0(n248), .A1(A[24]), .A2(n294), .B0(A[25]), .B1(n247), .Y(
        n292) );
  OAI32X1 U220 ( .A0(n246), .A1(A[26]), .A2(n295), .B0(A[27]), .B1(n245), .Y(
        n291) );
  OAI22XL U221 ( .A0(n296), .A1(n297), .B0(n298), .B1(n296), .Y(n265) );
  NOR3X1 U222 ( .A(n299), .B(n300), .C(n301), .Y(n298) );
  OAI21XL U223 ( .A0(B[8]), .A1(n239), .B0(n302), .Y(n299) );
  OAI31XL U224 ( .A0(n303), .A1(n304), .A2(n305), .B0(n306), .Y(n297) );
  AO22X1 U225 ( .A0(n240), .A1(n307), .B0(n305), .B1(n240), .Y(n306) );
  AOI32X1 U226 ( .A0(B[4]), .A1(n242), .A2(n308), .B0(n241), .B1(B[5]), .Y(
        n307) );
  AO21X1 U227 ( .A0(n260), .A1(A[6]), .B0(n310), .Y(n305) );
  AOI221XL U228 ( .A0(B[1]), .A1(n243), .B0(n311), .B1(B[0]), .C0(n312), .Y(
        n304) );
  OAI221XL U229 ( .A0(B[4]), .A1(n242), .B0(n313), .B1(n312), .C0(n308), .Y(
        n303) );
  OR2X1 U230 ( .A(B[5]), .B(n241), .Y(n308) );
  AND2X1 U231 ( .A(A[3]), .B(n261), .Y(n314) );
  OAI21XL U232 ( .A0(n300), .A1(n315), .B0(n316), .Y(n296) );
  OAI22XL U233 ( .A0(n317), .A1(n233), .B0(n318), .B1(n317), .Y(n316) );
  OAI32X1 U234 ( .A0(n258), .A1(A[14]), .A2(n321), .B0(A[15]), .B1(n257), .Y(
        n317) );
  AO22X1 U235 ( .A0(n322), .A1(n323), .B0(n301), .B1(n322), .Y(n315) );
  OAI21XL U236 ( .A0(B[10]), .A1(n237), .B0(n324), .Y(n301) );
  AOI21X1 U237 ( .A0(n258), .A1(A[14]), .B0(n321), .Y(n318) );
  NOR2BX1 U238 ( .AN(A[15]), .B(B[15]), .Y(n321) );
  OR2X1 U239 ( .A(B[13]), .B(n234), .Y(n320) );
  AO21X1 U240 ( .A0(n256), .A1(A[16]), .B0(n280), .Y(n264) );
  AND2X1 U241 ( .A(A[17]), .B(n255), .Y(n280) );
  NAND3X1 U242 ( .A(n269), .B(n282), .C(n279), .Y(n263) );
  AOI21X1 U243 ( .A0(n254), .A1(A[18]), .B0(n281), .Y(n279) );
  NOR2BX1 U244 ( .AN(A[19]), .B(B[19]), .Y(n281) );
  AOI211X1 U245 ( .A0(n252), .A1(A[20]), .B0(n275), .C0(n232), .Y(n282) );
  AOI21X1 U246 ( .A0(n250), .A1(A[22]), .B0(n276), .Y(n274) );
  NOR2BX1 U247 ( .AN(A[23]), .B(B[23]), .Y(n276) );
  AOI211X1 U248 ( .A0(n248), .A1(A[24]), .B0(n294), .C0(n325), .Y(n269) );
  NAND2BX1 U249 ( .AN(n283), .B(n293), .Y(n325) );
  AOI21X1 U250 ( .A0(n246), .A1(A[26]), .B0(n295), .Y(n293) );
  NOR2BX1 U251 ( .AN(A[27]), .B(B[27]), .Y(n295) );
  OAI211X1 U252 ( .A0(B[28]), .A1(n230), .B0(n289), .C0(n287), .Y(n283) );
  AOI21X1 U253 ( .A0(n244), .A1(A[30]), .B0(n290), .Y(n287) );
  NOR2BX1 U254 ( .AN(B[31]), .B(A[31]), .Y(n290) );
  OR2X1 U255 ( .A(B[29]), .B(n229), .Y(n289) );
  NOR2BX1 U256 ( .AN(A[25]), .B(B[25]), .Y(n294) );
endmodule


module SingleCycleProcessor_DW_leftsh_0 ( A, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  wire   n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n234, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361;

  MX2XL U178 ( .A(A[3]), .B(A[2]), .S0(n219), .Y(n350) );
  MX2XL U179 ( .A(A[21]), .B(A[20]), .S0(n218), .Y(n306) );
  MX2XL U180 ( .A(A[22]), .B(A[21]), .S0(n218), .Y(n302) );
  MX2XL U181 ( .A(A[1]), .B(A[0]), .S0(n219), .Y(n349) );
  MX2XL U182 ( .A(A[2]), .B(A[1]), .S0(n219), .Y(n356) );
  CLKINVX1 U183 ( .A(SH[2]), .Y(n224) );
  CLKINVX1 U184 ( .A(SH[3]), .Y(n225) );
  CLKINVX1 U185 ( .A(n308), .Y(n239) );
  CLKINVX1 U186 ( .A(n326), .Y(n243) );
  CLKINVX1 U187 ( .A(n299), .Y(n245) );
  CLKINVX1 U188 ( .A(n288), .Y(n234) );
  CLKINVX1 U189 ( .A(n318), .Y(n237) );
  CLKINVX1 U190 ( .A(n283), .Y(n242) );
  CLKINVX1 U191 ( .A(n251), .Y(n244) );
  CLKINVX1 U192 ( .A(n253), .Y(n246) );
  CLKINVX1 U193 ( .A(n256), .Y(n248) );
  CLKINVX1 U194 ( .A(n263), .Y(n230) );
  CLKINVX1 U195 ( .A(n307), .Y(B[22]) );
  CLKINVX1 U196 ( .A(n325), .Y(B[18]) );
  CLKINVX1 U197 ( .A(n335), .Y(B[16]) );
  CLKINVX1 U198 ( .A(n255), .Y(n247) );
  CLKINVX1 U199 ( .A(n257), .Y(n249) );
  CLKINVX1 U200 ( .A(n320), .Y(n250) );
  CLKINVX1 U201 ( .A(n278), .Y(n241) );
  CLKINVX1 U202 ( .A(n280), .Y(n232) );
  CLKINVX1 U203 ( .A(n273), .Y(n240) );
  CLKINVX1 U204 ( .A(n275), .Y(n231) );
  NOR2BX1 U205 ( .AN(n217), .B(n287), .Y(B[10]) );
  CLKINVX1 U206 ( .A(n228), .Y(n217) );
  CLKBUFX3 U207 ( .A(n221), .Y(n218) );
  CLKBUFX3 U208 ( .A(n221), .Y(n219) );
  CLKBUFX3 U209 ( .A(n228), .Y(n227) );
  CLKBUFX3 U210 ( .A(n228), .Y(n226) );
  CLKINVX1 U211 ( .A(n223), .Y(n222) );
  CLKBUFX3 U212 ( .A(n221), .Y(n220) );
  CLKINVX1 U213 ( .A(n268), .Y(n229) );
  CLKINVX1 U214 ( .A(n260), .Y(n238) );
  CLKBUFX3 U215 ( .A(SH[1]), .Y(n223) );
  CLKBUFX3 U216 ( .A(SH[0]), .Y(n221) );
  CLKBUFX3 U217 ( .A(SH[4]), .Y(n228) );
  NOR2X1 U218 ( .A(n227), .B(n251), .Y(B[9]) );
  NOR2X1 U219 ( .A(n227), .B(n252), .Y(B[8]) );
  NOR2X1 U220 ( .A(n227), .B(n253), .Y(B[7]) );
  NOR2X1 U221 ( .A(n227), .B(n254), .Y(B[6]) );
  NOR2X1 U222 ( .A(n227), .B(n255), .Y(B[5]) );
  NOR2X1 U223 ( .A(n227), .B(n256), .Y(B[4]) );
  NOR2X1 U224 ( .A(n227), .B(n257), .Y(B[3]) );
  MX3XL U225 ( .A(n258), .B(n259), .C(n238), .S0(SH[3]), .S1(n226), .Y(B[31])
         );
  MX3XL U226 ( .A(n261), .B(n262), .C(n230), .S0(n223), .S1(SH[2]), .Y(n258)
         );
  CLKMX2X2 U227 ( .A(A[31]), .B(A[30]), .S0(n219), .Y(n261) );
  MXI2X1 U228 ( .A(n264), .B(n265), .S0(n226), .Y(B[30]) );
  MX3XL U229 ( .A(n229), .B(n266), .C(n267), .S0(SH[2]), .S1(SH[3]), .Y(n264)
         );
  MX3XL U230 ( .A(A[30]), .B(A[29]), .C(n269), .S0(n220), .S1(n223), .Y(n268)
         );
  NOR2X1 U231 ( .A(n227), .B(n270), .Y(B[2]) );
  MX3XL U232 ( .A(n271), .B(n272), .C(n240), .S0(SH[3]), .S1(n227), .Y(B[29])
         );
  MX3XL U233 ( .A(n262), .B(n274), .C(n231), .S0(n223), .S1(SH[2]), .Y(n271)
         );
  CLKMX2X2 U234 ( .A(A[29]), .B(A[28]), .S0(n218), .Y(n262) );
  MX3XL U235 ( .A(n276), .B(n277), .C(n241), .S0(SH[3]), .S1(n227), .Y(B[28])
         );
  MX3XL U236 ( .A(n269), .B(n279), .C(n232), .S0(n223), .S1(SH[2]), .Y(n276)
         );
  CLKMX2X2 U237 ( .A(A[28]), .B(A[27]), .S0(n218), .Y(n269) );
  MX3XL U238 ( .A(n281), .B(n282), .C(n242), .S0(SH[3]), .S1(n226), .Y(B[27])
         );
  MXI2X1 U239 ( .A(n263), .B(n284), .S0(SH[2]), .Y(n281) );
  MXI2X1 U240 ( .A(n274), .B(n285), .S0(n223), .Y(n263) );
  CLKMX2X2 U241 ( .A(A[27]), .B(A[26]), .S0(n218), .Y(n274) );
  MXI2X1 U242 ( .A(n286), .B(n287), .S0(n226), .Y(B[26]) );
  MX3XL U243 ( .A(n266), .B(n288), .C(n289), .S0(SH[2]), .S1(SH[3]), .Y(n286)
         );
  MXI2X1 U244 ( .A(n279), .B(n290), .S0(n223), .Y(n266) );
  CLKMX2X2 U245 ( .A(A[26]), .B(A[25]), .S0(n218), .Y(n279) );
  MX3XL U246 ( .A(n291), .B(n292), .C(n244), .S0(SH[3]), .S1(n226), .Y(B[25])
         );
  MXI2X1 U247 ( .A(n293), .B(n294), .S0(SH[3]), .Y(n251) );
  MXI2X1 U248 ( .A(n275), .B(n295), .S0(SH[2]), .Y(n291) );
  MXI2X1 U249 ( .A(n285), .B(n296), .S0(n223), .Y(n275) );
  CLKMX2X2 U250 ( .A(A[25]), .B(A[24]), .S0(n218), .Y(n285) );
  MXI2X1 U251 ( .A(n297), .B(n252), .S0(n226), .Y(B[24]) );
  MXI2X1 U252 ( .A(n245), .B(n298), .S0(SH[3]), .Y(n252) );
  MX3XL U253 ( .A(n280), .B(n300), .C(n301), .S0(SH[2]), .S1(SH[3]), .Y(n297)
         );
  MXI2X1 U254 ( .A(n290), .B(n302), .S0(n223), .Y(n280) );
  CLKMX2X2 U255 ( .A(A[24]), .B(A[23]), .S0(n218), .Y(n290) );
  MX3XL U256 ( .A(n259), .B(n303), .C(n246), .S0(SH[3]), .S1(n226), .Y(B[23])
         );
  NAND2X1 U257 ( .A(n304), .B(n225), .Y(n253) );
  MXI2X1 U258 ( .A(n305), .B(n284), .S0(n224), .Y(n259) );
  MXI2X1 U259 ( .A(n296), .B(n306), .S0(n223), .Y(n284) );
  CLKMX2X2 U260 ( .A(A[23]), .B(A[22]), .S0(n218), .Y(n296) );
  MX3XL U261 ( .A(n267), .B(n308), .C(n254), .S0(SH[3]), .S1(n226), .Y(n307)
         );
  NAND2X1 U262 ( .A(n309), .B(n225), .Y(n254) );
  MXI2X1 U263 ( .A(n234), .B(n310), .S0(SH[2]), .Y(n267) );
  MXI2X1 U264 ( .A(n302), .B(n311), .S0(n223), .Y(n288) );
  MX3XL U265 ( .A(n272), .B(n312), .C(n247), .S0(SH[3]), .S1(n226), .Y(B[21])
         );
  NAND2X1 U266 ( .A(n313), .B(n225), .Y(n255) );
  MXI2X1 U267 ( .A(n314), .B(n295), .S0(n224), .Y(n272) );
  MXI2X1 U268 ( .A(n306), .B(n315), .S0(n223), .Y(n295) );
  MX3XL U269 ( .A(n277), .B(n316), .C(n248), .S0(SH[3]), .S1(n226), .Y(B[20])
         );
  NAND2X1 U270 ( .A(n317), .B(n225), .Y(n256) );
  MXI2X1 U271 ( .A(n318), .B(n300), .S0(n224), .Y(n277) );
  MXI2X1 U272 ( .A(n311), .B(n319), .S0(n223), .Y(n300) );
  CLKMX2X2 U273 ( .A(A[20]), .B(A[19]), .S0(n218), .Y(n311) );
  NOR2X1 U274 ( .A(n227), .B(n320), .Y(B[1]) );
  MX3XL U275 ( .A(n282), .B(n321), .C(n249), .S0(SH[3]), .S1(n226), .Y(B[19])
         );
  NAND2X1 U276 ( .A(n322), .B(n225), .Y(n257) );
  MXI2X1 U277 ( .A(n305), .B(n323), .S0(SH[2]), .Y(n282) );
  MXI2X1 U278 ( .A(n324), .B(n315), .S0(n222), .Y(n305) );
  CLKMX2X2 U279 ( .A(A[19]), .B(A[18]), .S0(n218), .Y(n315) );
  MX3XL U280 ( .A(n289), .B(n326), .C(n270), .S0(SH[3]), .S1(n226), .Y(n325)
         );
  NAND2X1 U281 ( .A(n327), .B(n225), .Y(n270) );
  MXI2X1 U282 ( .A(n310), .B(n328), .S0(SH[2]), .Y(n289) );
  CLKMX2X2 U283 ( .A(n329), .B(n319), .S0(n222), .Y(n310) );
  CLKMX2X2 U284 ( .A(A[18]), .B(A[17]), .S0(n218), .Y(n319) );
  MX3XL U285 ( .A(n292), .B(n293), .C(n250), .S0(SH[3]), .S1(n226), .Y(B[17])
         );
  NAND2X1 U286 ( .A(n294), .B(n225), .Y(n320) );
  NOR2X1 U287 ( .A(n330), .B(SH[2]), .Y(n294) );
  MXI2X1 U288 ( .A(n331), .B(n332), .S0(SH[2]), .Y(n293) );
  MXI2X1 U289 ( .A(n314), .B(n333), .S0(SH[2]), .Y(n292) );
  MXI2X1 U290 ( .A(n334), .B(n324), .S0(n222), .Y(n314) );
  CLKMX2X2 U291 ( .A(A[17]), .B(A[16]), .S0(n218), .Y(n324) );
  MX3XL U292 ( .A(n301), .B(n299), .C(n336), .S0(SH[3]), .S1(n226), .Y(n335)
         );
  MXI2X1 U293 ( .A(n337), .B(n338), .S0(n224), .Y(n299) );
  MXI2X1 U294 ( .A(n237), .B(n339), .S0(SH[2]), .Y(n301) );
  MXI2X1 U295 ( .A(n340), .B(n329), .S0(n222), .Y(n318) );
  CLKMX2X2 U296 ( .A(A[16]), .B(A[15]), .S0(n219), .Y(n329) );
  NOR2X1 U297 ( .A(n227), .B(n260), .Y(B[15]) );
  MXI2X1 U298 ( .A(n303), .B(n304), .S0(SH[3]), .Y(n260) );
  MXI2X1 U299 ( .A(n341), .B(n342), .S0(SH[2]), .Y(n304) );
  MXI2X1 U300 ( .A(n323), .B(n343), .S0(SH[2]), .Y(n303) );
  MXI2X1 U301 ( .A(n344), .B(n334), .S0(n222), .Y(n323) );
  CLKMX2X2 U302 ( .A(A[15]), .B(A[14]), .S0(n219), .Y(n334) );
  NOR2X1 U303 ( .A(n227), .B(n265), .Y(B[14]) );
  MXI2X1 U304 ( .A(n239), .B(n309), .S0(SH[3]), .Y(n265) );
  CLKMX2X2 U305 ( .A(n345), .B(n346), .S0(n224), .Y(n309) );
  MXI2X1 U306 ( .A(n347), .B(n328), .S0(n224), .Y(n308) );
  CLKMX2X2 U307 ( .A(n348), .B(n340), .S0(n222), .Y(n328) );
  CLKMX2X2 U308 ( .A(A[14]), .B(A[13]), .S0(n219), .Y(n340) );
  NOR2X1 U309 ( .A(n227), .B(n273), .Y(B[13]) );
  MXI2X1 U310 ( .A(n312), .B(n313), .S0(SH[3]), .Y(n273) );
  MXI2X1 U311 ( .A(n332), .B(n330), .S0(SH[2]), .Y(n313) );
  NAND2X1 U312 ( .A(n349), .B(n222), .Y(n330) );
  MXI2X1 U313 ( .A(n350), .B(n351), .S0(n222), .Y(n332) );
  MXI2X1 U314 ( .A(n333), .B(n331), .S0(SH[2]), .Y(n312) );
  MXI2X1 U315 ( .A(n352), .B(n353), .S0(n222), .Y(n331) );
  MXI2X1 U316 ( .A(n354), .B(n344), .S0(n222), .Y(n333) );
  CLKMX2X2 U317 ( .A(A[13]), .B(A[12]), .S0(n219), .Y(n344) );
  NOR2X1 U318 ( .A(n227), .B(n278), .Y(B[12]) );
  MXI2X1 U319 ( .A(n316), .B(n317), .S0(SH[3]), .Y(n278) );
  CLKMX2X2 U320 ( .A(n355), .B(n337), .S0(n224), .Y(n317) );
  CLKMX2X2 U321 ( .A(n356), .B(n357), .S0(n222), .Y(n337) );
  CLKMX2X2 U322 ( .A(n338), .B(n339), .S0(n224), .Y(n316) );
  CLKMX2X2 U323 ( .A(n358), .B(n348), .S0(n222), .Y(n339) );
  CLKMX2X2 U324 ( .A(A[12]), .B(A[11]), .S0(n219), .Y(n348) );
  CLKMX2X2 U325 ( .A(n359), .B(n360), .S0(n222), .Y(n338) );
  NOR2X1 U326 ( .A(n227), .B(n283), .Y(B[11]) );
  MXI2X1 U327 ( .A(n321), .B(n322), .S0(SH[3]), .Y(n283) );
  NOR2X1 U328 ( .A(n342), .B(SH[2]), .Y(n322) );
  MXI2X1 U329 ( .A(n350), .B(n349), .S0(n223), .Y(n342) );
  MXI2X1 U330 ( .A(n343), .B(n341), .S0(SH[2]), .Y(n321) );
  MXI2X1 U331 ( .A(n351), .B(n352), .S0(n222), .Y(n341) );
  CLKMX2X2 U332 ( .A(A[7]), .B(A[6]), .S0(n219), .Y(n352) );
  CLKMX2X2 U333 ( .A(A[5]), .B(A[4]), .S0(n219), .Y(n351) );
  MXI2X1 U334 ( .A(n353), .B(n354), .S0(n222), .Y(n343) );
  CLKMX2X2 U335 ( .A(A[11]), .B(A[10]), .S0(n219), .Y(n354) );
  CLKMX2X2 U336 ( .A(A[9]), .B(A[8]), .S0(n219), .Y(n353) );
  MXI2X1 U337 ( .A(n243), .B(n327), .S0(SH[3]), .Y(n287) );
  NOR2BX1 U338 ( .AN(n345), .B(SH[2]), .Y(n327) );
  CLKMX2X2 U339 ( .A(n361), .B(n356), .S0(n222), .Y(n345) );
  MXI2X1 U340 ( .A(n346), .B(n347), .S0(n224), .Y(n326) );
  CLKMX2X2 U341 ( .A(n360), .B(n358), .S0(n222), .Y(n347) );
  CLKMX2X2 U342 ( .A(A[10]), .B(A[9]), .S0(n220), .Y(n358) );
  CLKMX2X2 U343 ( .A(A[8]), .B(A[7]), .S0(n220), .Y(n360) );
  CLKMX2X2 U344 ( .A(n357), .B(n359), .S0(n222), .Y(n346) );
  CLKMX2X2 U345 ( .A(A[6]), .B(A[5]), .S0(n220), .Y(n359) );
  CLKMX2X2 U346 ( .A(A[4]), .B(A[3]), .S0(n220), .Y(n357) );
  NOR2X1 U347 ( .A(n227), .B(n336), .Y(B[0]) );
  NAND2X1 U348 ( .A(n298), .B(n225), .Y(n336) );
  NOR2BX1 U349 ( .AN(n355), .B(SH[2]), .Y(n298) );
  NOR2BX1 U350 ( .AN(n361), .B(n223), .Y(n355) );
  NOR2BX1 U351 ( .AN(A[0]), .B(n220), .Y(n361) );
endmodule


module SingleCycleProcessor_DW_rightsh_0 ( A, DATA_TC, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC;
  wire   n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366;

  INVXL U179 ( .A(A[2]), .Y(n253) );
  MX2XL U180 ( .A(A[2]), .B(A[3]), .S0(n221), .Y(n295) );
  MX2XL U181 ( .A(A[21]), .B(A[22]), .S0(n220), .Y(n342) );
  MX2XL U182 ( .A(A[20]), .B(A[21]), .S0(n221), .Y(n359) );
  MX2XL U183 ( .A(A[0]), .B(A[1]), .S0(n220), .Y(n366) );
  INVXL U184 ( .A(A[1]), .Y(n254) );
  CLKINVX1 U185 ( .A(SH[2]), .Y(n226) );
  CLKINVX1 U186 ( .A(SH[3]), .Y(n227) );
  CLKINVX1 U187 ( .A(n279), .Y(n239) );
  CLKINVX1 U188 ( .A(n285), .Y(n247) );
  CLKINVX1 U189 ( .A(n306), .Y(n244) );
  CLKINVX1 U190 ( .A(n310), .Y(n245) );
  CLKINVX1 U191 ( .A(n257), .Y(n246) );
  CLKINVX1 U192 ( .A(n275), .Y(n249) );
  CLKINVX1 U193 ( .A(n301), .Y(n231) );
  CLKINVX1 U194 ( .A(n291), .Y(n242) );
  CLKINVX1 U195 ( .A(n300), .Y(n238) );
  CLKINVX1 U196 ( .A(n302), .Y(n240) );
  CLKINVX1 U197 ( .A(n261), .Y(n237) );
  CLKINVX1 U198 ( .A(n332), .Y(n248) );
  CLKINVX1 U199 ( .A(n269), .Y(n243) );
  CLKINVX1 U200 ( .A(n280), .Y(n251) );
  CLKINVX1 U201 ( .A(n327), .Y(B[15]) );
  CLKINVX1 U202 ( .A(n338), .Y(B[13]) );
  CLKINVX1 U203 ( .A(n255), .Y(B[9]) );
  CLKINVX1 U204 ( .A(n270), .Y(n250) );
  CLKINVX1 U205 ( .A(n287), .Y(n252) );
  NOR2BX1 U206 ( .AN(n219), .B(n299), .Y(B[29]) );
  CLKINVX1 U207 ( .A(n230), .Y(n219) );
  CLKBUFX3 U208 ( .A(n223), .Y(n221) );
  CLKBUFX3 U209 ( .A(n223), .Y(n220) );
  CLKBUFX3 U210 ( .A(n230), .Y(n229) );
  CLKBUFX3 U211 ( .A(n230), .Y(n228) );
  CLKINVX1 U212 ( .A(n225), .Y(n224) );
  CLKBUFX3 U213 ( .A(n223), .Y(n222) );
  CLKINVX1 U214 ( .A(n326), .Y(n236) );
  CLKBUFX3 U215 ( .A(SH[1]), .Y(n225) );
  CLKBUFX3 U216 ( .A(SH[0]), .Y(n223) );
  CLKBUFX3 U217 ( .A(SH[4]), .Y(n230) );
  CLKINVX1 U218 ( .A(n282), .Y(B[3]) );
  CLKINVX1 U219 ( .A(n294), .Y(n241) );
  MX3XL U220 ( .A(n256), .B(n257), .C(n258), .S0(SH[3]), .S1(n228), .Y(n255)
         );
  MX3XL U221 ( .A(n259), .B(n260), .C(n237), .S0(SH[3]), .S1(n228), .Y(B[8])
         );
  MXI2X1 U222 ( .A(n262), .B(n263), .S0(n228), .Y(B[7]) );
  MX3XL U223 ( .A(n264), .B(n265), .C(n266), .S0(SH[2]), .S1(SH[3]), .Y(n262)
         );
  MX3XL U224 ( .A(n267), .B(n268), .C(n243), .S0(SH[3]), .S1(n228), .Y(B[6])
         );
  MXI2X1 U225 ( .A(n270), .B(n271), .S0(SH[2]), .Y(n267) );
  MXI2X1 U226 ( .A(n272), .B(n273), .S0(n228), .Y(B[5]) );
  MX3XL U227 ( .A(n274), .B(n275), .C(n276), .S0(SH[2]), .S1(SH[3]), .Y(n272)
         );
  MX3XL U228 ( .A(n277), .B(n278), .C(n239), .S0(SH[3]), .S1(n228), .Y(B[4])
         );
  MXI2X1 U229 ( .A(n280), .B(n281), .S0(SH[2]), .Y(n277) );
  MX3XL U230 ( .A(n283), .B(n247), .C(n284), .S0(SH[3]), .S1(n228), .Y(n282)
         );
  MX3XL U231 ( .A(n286), .B(n287), .C(n264), .S0(n225), .S1(SH[2]), .Y(n283)
         );
  MXI2X1 U232 ( .A(n288), .B(n289), .S0(n225), .Y(n264) );
  NOR2X1 U233 ( .A(n229), .B(n290), .Y(B[31]) );
  NOR2X1 U234 ( .A(n229), .B(n291), .Y(B[30]) );
  MX3XL U235 ( .A(n292), .B(n293), .C(n241), .S0(SH[3]), .S1(n228), .Y(B[2])
         );
  MX3XL U236 ( .A(n295), .B(n296), .C(n250), .S0(n225), .S1(SH[2]), .Y(n292)
         );
  MXI2X1 U237 ( .A(n297), .B(n298), .S0(n225), .Y(n270) );
  NOR2X1 U238 ( .A(n229), .B(n300), .Y(B[28]) );
  NOR2X1 U239 ( .A(n229), .B(n301), .Y(B[27]) );
  NOR2X1 U240 ( .A(n229), .B(n302), .Y(B[26]) );
  NOR2X1 U241 ( .A(n229), .B(n258), .Y(B[25]) );
  NAND2X1 U242 ( .A(n303), .B(n227), .Y(n258) );
  NOR2X1 U243 ( .A(n229), .B(n261), .Y(B[24]) );
  NAND2X1 U244 ( .A(n304), .B(n227), .Y(n261) );
  NOR2X1 U245 ( .A(n229), .B(n263), .Y(B[23]) );
  MXI2X1 U246 ( .A(n244), .B(n305), .S0(SH[3]), .Y(n263) );
  NOR2X1 U247 ( .A(n229), .B(n269), .Y(B[22]) );
  MXI2X1 U248 ( .A(n307), .B(n308), .S0(SH[3]), .Y(n269) );
  NOR2X1 U249 ( .A(n229), .B(n273), .Y(B[21]) );
  MXI2X1 U250 ( .A(n245), .B(n309), .S0(SH[3]), .Y(n273) );
  NOR2X1 U251 ( .A(n229), .B(n279), .Y(B[20]) );
  MXI2X1 U252 ( .A(n311), .B(n312), .S0(SH[3]), .Y(n279) );
  MXI2X1 U253 ( .A(n313), .B(n314), .S0(n228), .Y(B[1]) );
  MX3XL U254 ( .A(n315), .B(n274), .C(n256), .S0(SH[2]), .S1(SH[3]), .Y(n313)
         );
  MXI2X1 U255 ( .A(n249), .B(n316), .S0(SH[2]), .Y(n256) );
  MXI2X1 U256 ( .A(n289), .B(n317), .S0(n225), .Y(n275) );
  CLKMX2X2 U257 ( .A(A[9]), .B(A[10]), .S0(n221), .Y(n289) );
  MXI2X1 U258 ( .A(n252), .B(n288), .S0(n225), .Y(n274) );
  CLKMX2X2 U259 ( .A(A[7]), .B(A[8]), .S0(n220), .Y(n288) );
  MXI2X1 U260 ( .A(A[5]), .B(A[6]), .S0(n222), .Y(n287) );
  MX3XL U261 ( .A(n254), .B(n253), .C(n286), .S0(n222), .S1(n225), .Y(n315) );
  MXI2X1 U262 ( .A(A[3]), .B(A[4]), .S0(n222), .Y(n286) );
  NOR2X1 U263 ( .A(n229), .B(n284), .Y(B[19]) );
  MXI2X1 U264 ( .A(n318), .B(n319), .S0(SH[3]), .Y(n284) );
  NOR2X1 U265 ( .A(n229), .B(n294), .Y(B[18]) );
  MXI2X1 U266 ( .A(n320), .B(n321), .S0(SH[3]), .Y(n294) );
  NOR2X1 U267 ( .A(n229), .B(n314), .Y(B[17]) );
  MXI2X1 U268 ( .A(n246), .B(n303), .S0(SH[3]), .Y(n314) );
  CLKMX2X2 U269 ( .A(n322), .B(n323), .S0(n226), .Y(n303) );
  MXI2X1 U270 ( .A(n324), .B(n325), .S0(n226), .Y(n257) );
  NOR2X1 U271 ( .A(n229), .B(n326), .Y(B[16]) );
  MX3XL U272 ( .A(n266), .B(n306), .C(n290), .S0(SH[3]), .S1(n228), .Y(n327)
         );
  NAND2X1 U273 ( .A(n305), .B(n227), .Y(n290) );
  NOR2BX1 U274 ( .AN(n328), .B(SH[2]), .Y(n305) );
  MXI2X1 U275 ( .A(n329), .B(n330), .S0(n226), .Y(n306) );
  MXI2X1 U276 ( .A(n248), .B(n331), .S0(SH[2]), .Y(n266) );
  MX3XL U277 ( .A(n268), .B(n307), .C(n242), .S0(SH[3]), .S1(n228), .Y(B[14])
         );
  NAND2X1 U278 ( .A(n308), .B(n227), .Y(n291) );
  NOR2X1 U279 ( .A(n333), .B(SH[2]), .Y(n308) );
  MXI2X1 U280 ( .A(n334), .B(n335), .S0(SH[2]), .Y(n307) );
  MXI2X1 U281 ( .A(n336), .B(n337), .S0(SH[2]), .Y(n268) );
  MX3XL U282 ( .A(n276), .B(n310), .C(n299), .S0(SH[3]), .S1(n228), .Y(n338)
         );
  NAND2X1 U283 ( .A(n309), .B(n227), .Y(n299) );
  NOR2BX1 U284 ( .AN(n322), .B(SH[2]), .Y(n309) );
  CLKMX2X2 U285 ( .A(n339), .B(n340), .S0(n224), .Y(n322) );
  MXI2X1 U286 ( .A(n323), .B(n324), .S0(n226), .Y(n310) );
  CLKMX2X2 U287 ( .A(n341), .B(n342), .S0(n224), .Y(n324) );
  CLKMX2X2 U288 ( .A(n343), .B(n344), .S0(n224), .Y(n323) );
  MXI2X1 U289 ( .A(n316), .B(n325), .S0(SH[2]), .Y(n276) );
  CLKMX2X2 U290 ( .A(n345), .B(n346), .S0(n224), .Y(n325) );
  CLKMX2X2 U291 ( .A(n347), .B(n348), .S0(n224), .Y(n316) );
  MX3XL U292 ( .A(n278), .B(n311), .C(n238), .S0(SH[3]), .S1(n229), .Y(B[12])
         );
  NAND2X1 U293 ( .A(n312), .B(n227), .Y(n300) );
  NOR2X1 U294 ( .A(n349), .B(SH[2]), .Y(n312) );
  MXI2X1 U295 ( .A(n350), .B(n351), .S0(SH[2]), .Y(n311) );
  MXI2X1 U296 ( .A(n352), .B(n353), .S0(SH[2]), .Y(n278) );
  MX3XL U297 ( .A(n285), .B(n318), .C(n231), .S0(SH[3]), .S1(n229), .Y(B[11])
         );
  NAND2X1 U298 ( .A(n319), .B(n227), .Y(n301) );
  CLKMX2X2 U299 ( .A(n328), .B(n329), .S0(n226), .Y(n319) );
  CLKMX2X2 U300 ( .A(n340), .B(n343), .S0(n224), .Y(n329) );
  CLKMX2X2 U301 ( .A(A[27]), .B(A[28]), .S0(n220), .Y(n343) );
  CLKMX2X2 U302 ( .A(A[29]), .B(A[30]), .S0(n220), .Y(n340) );
  NOR2BX1 U303 ( .AN(n339), .B(n225), .Y(n328) );
  NOR2BX1 U304 ( .AN(A[31]), .B(n222), .Y(n339) );
  CLKMX2X2 U305 ( .A(n330), .B(n331), .S0(n226), .Y(n318) );
  CLKMX2X2 U306 ( .A(n342), .B(n345), .S0(n224), .Y(n331) );
  CLKMX2X2 U307 ( .A(A[19]), .B(A[20]), .S0(n220), .Y(n345) );
  CLKMX2X2 U308 ( .A(n344), .B(n341), .S0(n224), .Y(n330) );
  CLKMX2X2 U309 ( .A(A[23]), .B(A[24]), .S0(n220), .Y(n341) );
  CLKMX2X2 U310 ( .A(A[25]), .B(A[26]), .S0(n220), .Y(n344) );
  MXI2X1 U311 ( .A(n332), .B(n265), .S0(n226), .Y(n285) );
  MXI2X1 U312 ( .A(n317), .B(n348), .S0(n225), .Y(n265) );
  CLKMX2X2 U313 ( .A(A[13]), .B(A[14]), .S0(n220), .Y(n348) );
  CLKMX2X2 U314 ( .A(A[11]), .B(A[12]), .S0(n220), .Y(n317) );
  MXI2X1 U315 ( .A(n346), .B(n347), .S0(n224), .Y(n332) );
  CLKMX2X2 U316 ( .A(A[15]), .B(A[16]), .S0(n220), .Y(n347) );
  CLKMX2X2 U317 ( .A(A[17]), .B(A[18]), .S0(n220), .Y(n346) );
  MX3XL U318 ( .A(n293), .B(n320), .C(n240), .S0(SH[3]), .S1(n228), .Y(B[10])
         );
  NAND2X1 U319 ( .A(n321), .B(n227), .Y(n302) );
  MXI2X1 U320 ( .A(n335), .B(n333), .S0(SH[2]), .Y(n321) );
  NAND2X1 U321 ( .A(n354), .B(n224), .Y(n333) );
  MXI2X1 U322 ( .A(n355), .B(n356), .S0(n224), .Y(n335) );
  MXI2X1 U323 ( .A(n337), .B(n334), .S0(SH[2]), .Y(n320) );
  MXI2X1 U324 ( .A(n357), .B(n358), .S0(n224), .Y(n334) );
  MXI2X1 U325 ( .A(n359), .B(n360), .S0(n224), .Y(n337) );
  MXI2X1 U326 ( .A(n336), .B(n271), .S0(n226), .Y(n293) );
  MXI2X1 U327 ( .A(n361), .B(n362), .S0(n225), .Y(n271) );
  MXI2X1 U328 ( .A(n363), .B(n364), .S0(n224), .Y(n336) );
  MX3XL U329 ( .A(n365), .B(n259), .C(n236), .S0(SH[3]), .S1(n228), .Y(B[0])
         );
  MXI2X1 U330 ( .A(n260), .B(n304), .S0(SH[3]), .Y(n326) );
  MXI2X1 U331 ( .A(n351), .B(n349), .S0(SH[2]), .Y(n304) );
  MXI2X1 U332 ( .A(n355), .B(n354), .S0(n225), .Y(n349) );
  CLKMX2X2 U333 ( .A(A[30]), .B(A[31]), .S0(n220), .Y(n354) );
  CLKMX2X2 U334 ( .A(A[28]), .B(A[29]), .S0(n221), .Y(n355) );
  MXI2X1 U335 ( .A(n356), .B(n357), .S0(n224), .Y(n351) );
  CLKMX2X2 U336 ( .A(A[24]), .B(A[25]), .S0(n221), .Y(n357) );
  CLKMX2X2 U337 ( .A(A[26]), .B(A[27]), .S0(n221), .Y(n356) );
  MXI2X1 U338 ( .A(n353), .B(n350), .S0(SH[2]), .Y(n260) );
  MXI2X1 U339 ( .A(n358), .B(n359), .S0(n224), .Y(n350) );
  CLKMX2X2 U340 ( .A(A[22]), .B(A[23]), .S0(n221), .Y(n358) );
  MXI2X1 U341 ( .A(n360), .B(n363), .S0(n224), .Y(n353) );
  CLKMX2X2 U342 ( .A(A[16]), .B(A[17]), .S0(n221), .Y(n363) );
  CLKMX2X2 U343 ( .A(A[18]), .B(A[19]), .S0(n221), .Y(n360) );
  MXI2X1 U344 ( .A(n352), .B(n281), .S0(n226), .Y(n259) );
  MXI2X1 U345 ( .A(n298), .B(n361), .S0(n225), .Y(n281) );
  CLKMX2X2 U346 ( .A(A[10]), .B(A[11]), .S0(n221), .Y(n361) );
  CLKMX2X2 U347 ( .A(A[8]), .B(A[9]), .S0(n221), .Y(n298) );
  MXI2X1 U348 ( .A(n364), .B(n362), .S0(n224), .Y(n352) );
  CLKMX2X2 U349 ( .A(A[12]), .B(A[13]), .S0(n221), .Y(n362) );
  CLKMX2X2 U350 ( .A(A[14]), .B(A[15]), .S0(n221), .Y(n364) );
  MX3XL U351 ( .A(n366), .B(n295), .C(n251), .S0(n225), .S1(SH[2]), .Y(n365)
         );
  MXI2X1 U352 ( .A(n296), .B(n297), .S0(n225), .Y(n280) );
  CLKMX2X2 U353 ( .A(A[6]), .B(A[7]), .S0(n222), .Y(n297) );
  CLKMX2X2 U354 ( .A(A[4]), .B(A[5]), .S0(n222), .Y(n296) );
endmodule


module SingleCycleProcessor_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [31:1] carry;

  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX4 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  OR2X2 U1 ( .A(A[21]), .B(carry[21]), .Y(carry[22]) );
  XNOR2XL U2 ( .A(A[30]), .B(carry[30]), .Y(SUM[30]) );
  OR2X4 U3 ( .A(A[25]), .B(carry[25]), .Y(carry[26]) );
  OR2X4 U4 ( .A(A[23]), .B(carry[23]), .Y(carry[24]) );
  OR2X4 U5 ( .A(A[28]), .B(carry[28]), .Y(carry[29]) );
  OR2X4 U6 ( .A(A[17]), .B(carry[17]), .Y(carry[18]) );
  OR2X4 U7 ( .A(A[19]), .B(carry[19]), .Y(carry[20]) );
  XNOR2XL U8 ( .A(A[29]), .B(carry[29]), .Y(SUM[29]) );
  XNOR2XL U9 ( .A(A[28]), .B(carry[28]), .Y(SUM[28]) );
  XNOR2XL U10 ( .A(A[27]), .B(carry[27]), .Y(SUM[27]) );
  XNOR2XL U11 ( .A(A[26]), .B(carry[26]), .Y(SUM[26]) );
  XNOR2XL U12 ( .A(A[25]), .B(carry[25]), .Y(SUM[25]) );
  XNOR2XL U13 ( .A(A[24]), .B(carry[24]), .Y(SUM[24]) );
  INVXL U14 ( .A(A[0]), .Y(n4) );
  XNOR2XL U15 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XNOR2X1 U16 ( .A(A[31]), .B(carry[31]), .Y(SUM[31]) );
  NAND2X1 U17 ( .A(n1), .B(n2), .Y(carry[31]) );
  CLKINVX1 U18 ( .A(A[30]), .Y(n1) );
  CLKINVX1 U19 ( .A(carry[30]), .Y(n2) );
  OR2X1 U20 ( .A(A[15]), .B(carry[15]), .Y(carry[16]) );
  OR2X1 U21 ( .A(A[16]), .B(carry[16]), .Y(carry[17]) );
  OR2X1 U22 ( .A(A[18]), .B(carry[18]), .Y(carry[19]) );
  OR2X1 U23 ( .A(A[20]), .B(carry[20]), .Y(carry[21]) );
  OR2X1 U24 ( .A(A[29]), .B(carry[29]), .Y(carry[30]) );
  OR2X1 U25 ( .A(A[22]), .B(carry[22]), .Y(carry[23]) );
  OR2X1 U26 ( .A(A[24]), .B(carry[24]), .Y(carry[25]) );
  OR2X1 U27 ( .A(A[26]), .B(carry[26]), .Y(carry[27]) );
  OR2X1 U28 ( .A(A[27]), .B(carry[27]), .Y(carry[28]) );
  XNOR2XL U29 ( .A(A[15]), .B(carry[15]), .Y(SUM[15]) );
  XNOR2XL U30 ( .A(A[23]), .B(carry[23]), .Y(SUM[23]) );
  XNOR2XL U31 ( .A(A[22]), .B(carry[22]), .Y(SUM[22]) );
  XNOR2XL U32 ( .A(A[21]), .B(carry[21]), .Y(SUM[21]) );
  XNOR2XL U33 ( .A(A[20]), .B(carry[20]), .Y(SUM[20]) );
  XNOR2XL U34 ( .A(A[19]), .B(carry[19]), .Y(SUM[19]) );
  XNOR2XL U35 ( .A(A[18]), .B(carry[18]), .Y(SUM[18]) );
  XNOR2XL U36 ( .A(A[17]), .B(carry[17]), .Y(SUM[17]) );
  XNOR2XL U37 ( .A(A[16]), .B(carry[16]), .Y(SUM[16]) );
  NAND2X1 U38 ( .A(n3), .B(n4), .Y(carry[1]) );
  CLKINVX1 U39 ( .A(B[0]), .Y(n3) );
endmodule


module SingleCycleProcessor_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20;
  wire   [31:1] carry;

  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  CLKINVX4 U1 ( .A(A[0]), .Y(n19) );
  NAND2BX1 U2 ( .AN(n15), .B(A[29]), .Y(n16) );
  OR2X1 U3 ( .A(n16), .B(n17), .Y(n1) );
  NAND2BX1 U4 ( .AN(n14), .B(A[28]), .Y(n15) );
  NAND2BX1 U5 ( .AN(n13), .B(A[27]), .Y(n14) );
  NAND2BX1 U6 ( .AN(n9), .B(A[23]), .Y(n10) );
  NAND2BX1 U7 ( .AN(n5), .B(A[19]), .Y(n6) );
  NAND2BX1 U8 ( .AN(n7), .B(A[21]), .Y(n8) );
  NAND2BX1 U9 ( .AN(n11), .B(A[25]), .Y(n12) );
  NAND2BX1 U10 ( .AN(n3), .B(A[17]), .Y(n4) );
  NAND2BX1 U11 ( .AN(n18), .B(A[15]), .Y(n2) );
  XNOR2X1 U12 ( .A(A[31]), .B(n1), .Y(SUM[31]) );
  CLKINVX1 U13 ( .A(A[30]), .Y(n17) );
  NOR2XL U14 ( .A(n19), .B(n20), .Y(carry[1]) );
  XNOR2XL U15 ( .A(B[0]), .B(n19), .Y(SUM[0]) );
  CLKINVX1 U16 ( .A(carry[15]), .Y(n18) );
  XNOR2XL U17 ( .A(A[30]), .B(n16), .Y(SUM[30]) );
  XNOR2X1 U18 ( .A(A[29]), .B(n15), .Y(SUM[29]) );
  XNOR2X1 U19 ( .A(A[28]), .B(n14), .Y(SUM[28]) );
  XNOR2X1 U20 ( .A(A[27]), .B(n13), .Y(SUM[27]) );
  XNOR2XL U21 ( .A(A[26]), .B(n12), .Y(SUM[26]) );
  XNOR2X1 U22 ( .A(A[25]), .B(n11), .Y(SUM[25]) );
  CLKINVX1 U23 ( .A(B[0]), .Y(n20) );
  NAND2BX1 U24 ( .AN(n2), .B(A[16]), .Y(n3) );
  NAND2BX1 U25 ( .AN(n4), .B(A[18]), .Y(n5) );
  NAND2BX1 U26 ( .AN(n6), .B(A[20]), .Y(n7) );
  NAND2BX1 U27 ( .AN(n8), .B(A[22]), .Y(n9) );
  NAND2BX1 U28 ( .AN(n10), .B(A[24]), .Y(n11) );
  NAND2BX1 U29 ( .AN(n12), .B(A[26]), .Y(n13) );
  XNOR2XL U30 ( .A(A[24]), .B(n10), .Y(SUM[24]) );
  XNOR2XL U31 ( .A(A[23]), .B(n9), .Y(SUM[23]) );
  XNOR2XL U32 ( .A(A[22]), .B(n8), .Y(SUM[22]) );
  XNOR2XL U33 ( .A(A[21]), .B(n7), .Y(SUM[21]) );
  XNOR2XL U34 ( .A(A[20]), .B(n6), .Y(SUM[20]) );
  XNOR2XL U35 ( .A(A[19]), .B(n5), .Y(SUM[19]) );
  XNOR2XL U36 ( .A(A[18]), .B(n4), .Y(SUM[18]) );
  XNOR2XL U37 ( .A(A[17]), .B(n3), .Y(SUM[17]) );
  XNOR2XL U38 ( .A(A[16]), .B(n2), .Y(SUM[16]) );
  XNOR2XL U39 ( .A(A[15]), .B(n18), .Y(SUM[15]) );
endmodule


module SingleCycleProcessor_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \carry[31] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26;
  wire   [31:1] carry;

  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(\carry[28] ), .CO(\carry[29] ), .S(
        SUM[28]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(\carry[25] ), .CO(\carry[26] ), .S(
        SUM[25]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(\carry[18] ), .CO(\carry[19] ), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(\carry[17] ), .CO(\carry[18] ), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(\carry[16] ), .CO(\carry[17] ), .S(
        SUM[16]) );
  ADDFHX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(\carry[29] ), .CO(\carry[30] ), 
        .S(SUM[29]) );
  ADDFHX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(\carry[26] ), .CO(\carry[27] ), 
        .S(SUM[26]) );
  ADDFHX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(\carry[27] ), .CO(\carry[28] ), 
        .S(SUM[27]) );
  ADDFHX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX4 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX4 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(\carry[30] ), .CO(\carry[31] ), .S(
        SUM[30]) );
  ADDFHX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(\carry[23] ), .CO(\carry[24] ), 
        .S(SUM[23]) );
  ADDFHX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(\carry[24] ), .CO(\carry[25] ), 
        .S(SUM[24]) );
  ADDFHX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(\carry[22] ), .CO(\carry[23] ), 
        .S(SUM[22]) );
  CMPR32X2 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .CO(\carry[15] ), .S(
        SUM[14]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(\carry[21] ), .CO(\carry[22] ), .S(
        SUM[21]) );
  ADDFHX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(\carry[19] ), .CO(\carry[20] ), 
        .S(SUM[19]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(\carry[20] ), .CO(\carry[21] ), .S(
        SUM[20]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(\carry[15] ), .CO(\carry[16] ), .S(
        SUM[15]) );
  CLKINVX2 U1 ( .A(A[0]), .Y(n25) );
  NAND2XL U2 ( .A(carry[1]), .B(A[1]), .Y(n18) );
  NAND2XL U3 ( .A(B[1]), .B(A[1]), .Y(n19) );
  NAND2X1 U4 ( .A(B[1]), .B(carry[1]), .Y(n20) );
  NAND2XL U5 ( .A(B[4]), .B(A[4]), .Y(n5) );
  NAND2XL U6 ( .A(A[4]), .B(carry[4]), .Y(n3) );
  NAND2X1 U7 ( .A(B[12]), .B(A[12]), .Y(n12) );
  NAND2X2 U8 ( .A(B[12]), .B(carry[12]), .Y(n11) );
  NOR2X1 U9 ( .A(n25), .B(n26), .Y(carry[1]) );
  NAND2X2 U10 ( .A(B[2]), .B(A[2]), .Y(n24) );
  XOR2XL U11 ( .A(B[31]), .B(A[31]), .Y(n1) );
  XOR2X1 U12 ( .A(n1), .B(\carry[31] ), .Y(SUM[31]) );
  XOR2XL U13 ( .A(B[4]), .B(A[4]), .Y(n2) );
  XOR2XL U14 ( .A(n2), .B(carry[4]), .Y(SUM[4]) );
  NAND2X2 U15 ( .A(B[4]), .B(carry[4]), .Y(n4) );
  NAND3X2 U16 ( .A(n3), .B(n4), .C(n5), .Y(carry[5]) );
  XOR2X1 U17 ( .A(B[6]), .B(A[6]), .Y(n6) );
  XOR2XL U18 ( .A(n6), .B(carry[6]), .Y(SUM[6]) );
  NAND2X2 U19 ( .A(A[6]), .B(carry[6]), .Y(n7) );
  NAND2X2 U20 ( .A(B[6]), .B(carry[6]), .Y(n8) );
  NAND2X2 U21 ( .A(B[6]), .B(A[6]), .Y(n9) );
  NAND3X2 U22 ( .A(n7), .B(n8), .C(n9), .Y(carry[7]) );
  XOR3XL U23 ( .A(carry[12]), .B(B[12]), .C(A[12]), .Y(SUM[12]) );
  NAND2X2 U24 ( .A(A[12]), .B(carry[12]), .Y(n10) );
  NAND3X2 U25 ( .A(n10), .B(n11), .C(n12), .Y(carry[13]) );
  XOR2XL U26 ( .A(B[10]), .B(A[10]), .Y(n13) );
  XOR2XL U27 ( .A(n13), .B(carry[10]), .Y(SUM[10]) );
  NAND2X2 U28 ( .A(A[10]), .B(carry[10]), .Y(n14) );
  NAND2X2 U29 ( .A(B[10]), .B(carry[10]), .Y(n15) );
  NAND2X2 U30 ( .A(B[10]), .B(A[10]), .Y(n16) );
  NAND3X2 U31 ( .A(n14), .B(n15), .C(n16), .Y(carry[11]) );
  XOR2XL U32 ( .A(B[1]), .B(carry[1]), .Y(n17) );
  XOR2XL U33 ( .A(n17), .B(A[1]), .Y(SUM[1]) );
  NAND3X2 U34 ( .A(n18), .B(n19), .C(n20), .Y(carry[2]) );
  NAND2X1 U35 ( .A(A[2]), .B(carry[2]), .Y(n22) );
  NAND2X1 U36 ( .A(B[2]), .B(carry[2]), .Y(n23) );
  NAND3X1 U37 ( .A(n22), .B(n23), .C(n24), .Y(carry[3]) );
  XOR2XL U38 ( .A(B[2]), .B(A[2]), .Y(n21) );
  XOR2XL U39 ( .A(n21), .B(carry[2]), .Y(SUM[2]) );
  XNOR2XL U40 ( .A(B[0]), .B(n25), .Y(SUM[0]) );
  CLKINVX1 U41 ( .A(B[0]), .Y(n26) );
endmodule


module SingleCycleProcessor_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50;
  wire   [32:0] carry;

  ADDFXL U2_4 ( .A(A[4]), .B(n46), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_27 ( .A(A[27]), .B(n23), .CI(carry[27]), .CO(carry[28]), .S(
        DIFF[27]) );
  ADDFXL U2_25 ( .A(A[25]), .B(n25), .CI(carry[25]), .CO(carry[26]), .S(
        DIFF[25]) );
  ADDFXL U2_7 ( .A(A[7]), .B(n43), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n45), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFHX1 U2_6 ( .A(A[6]), .B(n44), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFHX1 U2_26 ( .A(A[26]), .B(n24), .CI(carry[26]), .CO(carry[27]), .S(
        DIFF[26]) );
  ADDFHX2 U2_24 ( .A(A[24]), .B(n26), .CI(carry[24]), .CO(carry[25]), .S(
        DIFF[24]) );
  ADDFHX2 U2_18 ( .A(A[18]), .B(n32), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  ADDFHX2 U2_14 ( .A(A[14]), .B(n36), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFHX1 U2_8 ( .A(A[8]), .B(n42), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8])
         );
  ADDFHX1 U2_29 ( .A(A[29]), .B(n21), .CI(carry[29]), .CO(carry[30]), .S(
        DIFF[29]) );
  ADDFHX2 U2_9 ( .A(A[9]), .B(n41), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFHX1 U2_28 ( .A(A[28]), .B(n22), .CI(carry[28]), .CO(carry[29]), .S(
        DIFF[28]) );
  ADDFHX1 U2_1 ( .A(A[1]), .B(n49), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  ADDFHX2 U2_13 ( .A(A[13]), .B(n37), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFHX2 U2_21 ( .A(A[21]), .B(n29), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  ADDFHX2 U2_16 ( .A(A[16]), .B(n34), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  ADDFX2 U2_17 ( .A(A[17]), .B(n33), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  ADDFHX2 U2_19 ( .A(A[19]), .B(n31), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  ADDFHX2 U2_22 ( .A(A[22]), .B(n28), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  ADDFHX2 U2_15 ( .A(A[15]), .B(n35), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  ADDFHX2 U2_20 ( .A(A[20]), .B(n30), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  ADDFHX2 U2_11 ( .A(A[11]), .B(n39), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_3 ( .A(A[3]), .B(n47), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFHX2 U2_30 ( .A(A[30]), .B(n20), .CI(carry[30]), .CO(carry[31]), .S(
        DIFF[30]) );
  XOR3X2 U2_31 ( .A(A[31]), .B(n19), .C(carry[31]), .Y(DIFF[31]) );
  INVXL U1 ( .A(A[0]), .Y(n18) );
  NAND2X1 U2 ( .A(A[23]), .B(carry[23]), .Y(n6) );
  NAND2X1 U3 ( .A(n27), .B(carry[23]), .Y(n7) );
  NAND2X1 U4 ( .A(n40), .B(A[10]), .Y(n16) );
  NAND2X1 U5 ( .A(n48), .B(carry[2]), .Y(n10) );
  NAND2X2 U6 ( .A(n38), .B(carry[12]), .Y(n3) );
  CLKINVX1 U7 ( .A(B[23]), .Y(n27) );
  NAND3X1 U8 ( .A(n10), .B(n11), .C(n12), .Y(carry[3]) );
  NAND2XL U9 ( .A(A[2]), .B(carry[2]), .Y(n11) );
  XOR2XL U10 ( .A(n38), .B(A[12]), .Y(n1) );
  XOR2XL U11 ( .A(n1), .B(carry[12]), .Y(DIFF[12]) );
  NAND2X2 U12 ( .A(A[12]), .B(carry[12]), .Y(n2) );
  NAND2X2 U13 ( .A(n38), .B(A[12]), .Y(n4) );
  NAND3X2 U14 ( .A(n2), .B(n3), .C(n4), .Y(carry[13]) );
  INVX1 U15 ( .A(B[12]), .Y(n38) );
  XOR2XL U16 ( .A(n27), .B(A[23]), .Y(n5) );
  XOR2XL U17 ( .A(n5), .B(carry[23]), .Y(DIFF[23]) );
  NAND2X4 U18 ( .A(n27), .B(A[23]), .Y(n8) );
  NAND3X2 U19 ( .A(n6), .B(n7), .C(n8), .Y(carry[24]) );
  XOR2XL U20 ( .A(A[2]), .B(n48), .Y(n9) );
  XOR2XL U21 ( .A(n9), .B(carry[2]), .Y(DIFF[2]) );
  NAND2XL U22 ( .A(A[2]), .B(n48), .Y(n12) );
  XOR2XL U23 ( .A(n40), .B(A[10]), .Y(n13) );
  XOR2XL U24 ( .A(n13), .B(carry[10]), .Y(DIFF[10]) );
  NAND2X2 U25 ( .A(A[10]), .B(carry[10]), .Y(n14) );
  NAND2X2 U26 ( .A(n40), .B(carry[10]), .Y(n15) );
  NAND3X2 U27 ( .A(n14), .B(n15), .C(n16), .Y(carry[11]) );
  CLKINVX1 U28 ( .A(B[10]), .Y(n40) );
  INVXL U29 ( .A(B[2]), .Y(n48) );
  INVXL U30 ( .A(B[0]), .Y(n50) );
  INVX1 U31 ( .A(B[1]), .Y(n49) );
  INVX1 U32 ( .A(B[3]), .Y(n47) );
  INVXL U33 ( .A(B[11]), .Y(n39) );
  INVXL U34 ( .A(B[9]), .Y(n41) );
  INVXL U35 ( .A(B[8]), .Y(n42) );
  INVXL U36 ( .A(B[6]), .Y(n44) );
  XNOR2XL U37 ( .A(n50), .B(A[0]), .Y(DIFF[0]) );
  NAND2X1 U38 ( .A(n17), .B(n18), .Y(carry[1]) );
  CLKINVX1 U39 ( .A(n50), .Y(n17) );
  CLKINVX1 U40 ( .A(B[5]), .Y(n45) );
  CLKINVX1 U41 ( .A(B[7]), .Y(n43) );
  CLKINVX1 U42 ( .A(B[13]), .Y(n37) );
  CLKINVX1 U43 ( .A(B[14]), .Y(n36) );
  CLKINVX1 U44 ( .A(B[15]), .Y(n35) );
  CLKINVX1 U45 ( .A(B[16]), .Y(n34) );
  CLKINVX1 U46 ( .A(B[17]), .Y(n33) );
  CLKINVX1 U47 ( .A(B[18]), .Y(n32) );
  CLKINVX1 U48 ( .A(B[19]), .Y(n31) );
  CLKINVX1 U49 ( .A(B[20]), .Y(n30) );
  CLKINVX1 U50 ( .A(B[21]), .Y(n29) );
  CLKINVX1 U51 ( .A(B[22]), .Y(n28) );
  CLKINVX1 U52 ( .A(B[24]), .Y(n26) );
  CLKINVX1 U53 ( .A(B[25]), .Y(n25) );
  CLKINVX1 U54 ( .A(B[26]), .Y(n24) );
  CLKINVX1 U55 ( .A(B[27]), .Y(n23) );
  CLKINVX1 U56 ( .A(B[28]), .Y(n22) );
  CLKINVX1 U57 ( .A(B[29]), .Y(n21) );
  CLKINVX1 U58 ( .A(B[30]), .Y(n20) );
  CLKINVX1 U59 ( .A(B[4]), .Y(n46) );
  CLKINVX1 U60 ( .A(B[31]), .Y(n19) );
endmodule


module SingleCycleProcessor_DW01_add_3 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  wire   [31:1] carry;

  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFHX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFHX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFHX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFHX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX4 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFHX4 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  INVXL U1 ( .A(A[0]), .Y(n9) );
  NAND2X1 U2 ( .A(A[14]), .B(carry[14]), .Y(n6) );
  NAND2X1 U3 ( .A(B[14]), .B(carry[14]), .Y(n7) );
  NAND2X1 U4 ( .A(B[14]), .B(A[14]), .Y(n8) );
  NAND3X1 U5 ( .A(n6), .B(n7), .C(n8), .Y(carry[15]) );
  XOR2XL U6 ( .A(A[3]), .B(B[3]), .Y(n1) );
  XOR2XL U7 ( .A(n1), .B(carry[3]), .Y(SUM[3]) );
  NAND2X1 U8 ( .A(B[3]), .B(carry[3]), .Y(n2) );
  NAND2X1 U9 ( .A(A[3]), .B(carry[3]), .Y(n3) );
  NAND2XL U10 ( .A(A[3]), .B(B[3]), .Y(n4) );
  NAND3X1 U11 ( .A(n2), .B(n3), .C(n4), .Y(carry[4]) );
  XOR2XL U12 ( .A(B[14]), .B(A[14]), .Y(n5) );
  XOR2XL U13 ( .A(n5), .B(carry[14]), .Y(SUM[14]) );
  NOR2XL U14 ( .A(n9), .B(n10), .Y(carry[1]) );
  XNOR2XL U15 ( .A(B[0]), .B(n9), .Y(SUM[0]) );
  CLKINVX1 U16 ( .A(B[0]), .Y(n10) );
endmodule


module SingleCycleProcessor_DW01_inc_0 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  ADDHXL U1_1_30 ( .A(A[30]), .B(carry[30]), .CO(carry[31]), .S(SUM[30]) );
  ADDHXL U1_1_29 ( .A(A[29]), .B(carry[29]), .CO(carry[30]), .S(SUM[29]) );
  ADDHXL U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  ADDHXL U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  ADDHXL U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  ADDHXL U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  ADDHXL U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  ADDHXL U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  ADDHXL U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  ADDHXL U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  ADDHXL U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  ADDHXL U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  ADDHXL U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  ADDHXL U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  ADDHXL U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  ADDHXL U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADDHXL U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXL U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[31]), .B(A[31]), .Y(SUM[31]) );
endmodule


module SingleCycleProcessor_DW01_add_4 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \carry[31] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , n1, n2;
  wire   [31:1] carry;

  XOR3X1 U1_31 ( .A(A[31]), .B(B[31]), .C(\carry[31] ), .Y(SUM[31]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(\carry[20] ), .CO(\carry[21] ), .S(
        SUM[20]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(\carry[18] ), .CO(\carry[19] ), .S(
        SUM[18]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(\carry[16] ), .CO(\carry[17] ), .S(
        SUM[16]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(\carry[25] ), .CO(\carry[26] ), 
        .S(SUM[25]) );
  ADDFHX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(\carry[19] ), .CO(\carry[20] ), 
        .S(SUM[19]) );
  ADDFHX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(\carry[17] ), .CO(\carry[18] ), 
        .S(SUM[17]) );
  ADDFHX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(\carry[28] ), .CO(\carry[29] ), 
        .S(SUM[28]) );
  ADDFHX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(\carry[22] ), .CO(\carry[23] ), 
        .S(SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(\carry[21] ), .CO(\carry[22] ), .S(
        SUM[21]) );
  ADDFHX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(\carry[15] ), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(\carry[15] ), .CO(\carry[16] ), .S(
        SUM[15]) );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(\carry[29] ), .CO(\carry[30] ), 
        .S(SUM[29]) );
  ADDFHX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(\carry[30] ), .CO(\carry[31] ), 
        .S(SUM[30]) );
  ADDFHX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(\carry[26] ), .CO(\carry[27] ), 
        .S(SUM[26]) );
  ADDFHX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(\carry[27] ), .CO(\carry[28] ), 
        .S(SUM[27]) );
  ADDFHX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(\carry[23] ), .CO(\carry[24] ), 
        .S(SUM[23]) );
  ADDFHX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(\carry[24] ), .CO(\carry[25] ), 
        .S(SUM[24]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(n2) );
  XNOR2XL U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND2X1 U3 ( .A(n1), .B(n2), .Y(carry[1]) );
  CLKINVX1 U4 ( .A(B[0]), .Y(n1) );
endmodule


module SingleCycleProcessor_DW01_inc_1 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  ADDHXL U1_1_30 ( .A(A[30]), .B(carry[30]), .CO(carry[31]), .S(SUM[30]) );
  ADDHXL U1_1_29 ( .A(A[29]), .B(carry[29]), .CO(carry[30]), .S(SUM[29]) );
  ADDHXL U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  ADDHXL U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  ADDHXL U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  ADDHXL U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  ADDHXL U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  ADDHXL U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  ADDHXL U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  ADDHXL U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  ADDHXL U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  ADDHXL U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  ADDHXL U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  ADDHXL U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  ADDHXL U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  ADDHXL U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADDHXL U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXL U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INVXL U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[31]), .B(A[31]), .Y(SUM[31]) );
endmodule


module SingleCycleProcessor_DW01_add_5 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;
  wire   [31:1] carry;

  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFHX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFHX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X2 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFHX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFHX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFHX4 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX4 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  NAND2X1 U1 ( .A(A[22]), .B(carry[22]), .Y(n7) );
  NAND3X1 U2 ( .A(n6), .B(n7), .C(n8), .Y(carry[23]) );
  NAND2X1 U3 ( .A(A[22]), .B(B[22]), .Y(n8) );
  NAND2X1 U4 ( .A(B[22]), .B(carry[22]), .Y(n6) );
  NAND2XL U5 ( .A(B[2]), .B(carry[2]), .Y(n2) );
  XOR2XL U6 ( .A(A[2]), .B(B[2]), .Y(n1) );
  XOR2XL U7 ( .A(n1), .B(carry[2]), .Y(SUM[2]) );
  NAND2X1 U8 ( .A(A[2]), .B(carry[2]), .Y(n3) );
  NAND2XL U9 ( .A(A[2]), .B(B[2]), .Y(n4) );
  NAND3X1 U10 ( .A(n2), .B(n3), .C(n4), .Y(carry[3]) );
  XOR2XL U11 ( .A(A[22]), .B(B[22]), .Y(n5) );
  XOR2XL U12 ( .A(n5), .B(carry[22]), .Y(SUM[22]) );
  XOR2XL U13 ( .A(A[6]), .B(B[6]), .Y(n9) );
  XOR2XL U14 ( .A(n9), .B(carry[6]), .Y(SUM[6]) );
  NAND2X2 U15 ( .A(B[6]), .B(carry[6]), .Y(n10) );
  NAND2X2 U16 ( .A(A[6]), .B(carry[6]), .Y(n11) );
  NAND2X2 U17 ( .A(A[6]), .B(B[6]), .Y(n12) );
  NAND3X2 U18 ( .A(n10), .B(n11), .C(n12), .Y(carry[7]) );
  XNOR2XL U19 ( .A(B[0]), .B(n13), .Y(SUM[0]) );
  CLKINVX1 U20 ( .A(A[0]), .Y(n13) );
  NOR2X1 U21 ( .A(n13), .B(n14), .Y(carry[1]) );
  CLKINVX1 U22 ( .A(B[0]), .Y(n14) );
endmodule


module SingleCycleProcessor ( PC, datain, address, MW, MR, instruction, 
        dataout, clk, reset_n );
  output [31:0] PC;
  output [31:0] datain;
  output [31:0] address;
  input [31:0] instruction;
  input [31:0] dataout;
  input clk, reset_n;
  output MW, MR;
  wire   N46, N47, N48, N49, N50, N51, N52, N53, N54, \R[1][31] , \R[1][30] ,
         \R[1][29] , \R[1][28] , \R[1][27] , \R[1][26] , \R[1][25] ,
         \R[1][24] , \R[1][23] , \R[1][22] , \R[1][21] , \R[1][20] ,
         \R[1][19] , \R[1][18] , \R[1][17] , \R[1][16] , \R[1][15] ,
         \R[1][14] , \R[1][13] , \R[1][12] , \R[1][11] , \R[1][10] , \R[1][9] ,
         \R[1][8] , \R[1][7] , \R[1][6] , \R[1][5] , \R[1][4] , \R[1][3] ,
         \R[1][2] , \R[1][1] , \R[1][0] , \R[3][31] , \R[3][30] , \R[3][29] ,
         \R[3][28] , \R[3][27] , \R[3][26] , \R[3][25] , \R[3][24] ,
         \R[3][23] , \R[3][22] , \R[3][21] , \R[3][20] , \R[3][19] ,
         \R[3][18] , \R[3][17] , \R[3][16] , \R[3][15] , \R[3][14] ,
         \R[3][13] , \R[3][12] , \R[3][11] , \R[3][10] , \R[3][9] , \R[3][8] ,
         \R[3][7] , \R[3][6] , \R[3][5] , \R[3][4] , \R[3][3] , \R[3][2] ,
         \R[3][1] , \R[3][0] , \R[4][31] , \R[4][30] , \R[4][29] , \R[4][28] ,
         \R[4][27] , \R[4][26] , \R[4][25] , \R[4][24] , \R[4][23] ,
         \R[4][22] , \R[4][21] , \R[4][20] , \R[4][19] , \R[4][18] ,
         \R[4][17] , \R[4][16] , \R[4][15] , \R[4][14] , \R[4][13] ,
         \R[4][12] , \R[4][11] , \R[4][10] , \R[4][9] , \R[4][8] , \R[4][7] ,
         \R[4][6] , \R[4][5] , \R[4][4] , \R[4][3] , \R[4][2] , \R[4][1] ,
         \R[4][0] , \R[5][31] , \R[5][30] , \R[5][29] , \R[5][28] , \R[5][27] ,
         \R[5][26] , \R[5][25] , \R[5][24] , \R[5][23] , \R[5][22] ,
         \R[5][21] , \R[5][20] , \R[5][19] , \R[5][18] , \R[5][17] ,
         \R[5][16] , \R[5][15] , \R[5][14] , \R[5][13] , \R[5][12] ,
         \R[5][11] , \R[5][10] , \R[5][9] , \R[5][8] , \R[5][7] , \R[5][6] ,
         \R[5][5] , \R[5][4] , \R[5][3] , \R[5][2] , \R[5][1] , \R[5][0] ,
         \R[6][31] , \R[6][30] , \R[6][29] , \R[6][28] , \R[6][27] ,
         \R[6][26] , \R[6][25] , \R[6][24] , \R[6][23] , \R[6][22] ,
         \R[6][21] , \R[6][20] , \R[6][19] , \R[6][18] , \R[6][17] ,
         \R[6][16] , \R[6][15] , \R[6][14] , \R[6][13] , \R[6][12] ,
         \R[6][11] , \R[6][10] , \R[6][9] , \R[6][8] , \R[6][7] , \R[6][6] ,
         \R[6][5] , \R[6][4] , \R[6][3] , \R[6][2] , \R[6][1] , \R[6][0] ,
         \R[7][31] , \R[7][30] , \R[7][29] , \R[7][28] , \R[7][27] ,
         \R[7][26] , \R[7][25] , \R[7][24] , \R[7][23] , \R[7][22] ,
         \R[7][21] , \R[7][20] , \R[7][19] , \R[7][18] , \R[7][17] ,
         \R[7][16] , \R[7][15] , \R[7][14] , \R[7][13] , \R[7][12] ,
         \R[7][11] , \R[7][10] , \R[7][9] , \R[7][8] , \R[7][7] , \R[7][6] ,
         \R[7][5] , \R[7][4] , \R[7][3] , \R[7][2] , \R[7][1] , \R[7][0] ,
         \R[8][31] , \R[8][30] , \R[8][29] , \R[8][28] , \R[8][27] ,
         \R[8][26] , \R[8][25] , \R[8][24] , \R[8][23] , \R[8][22] ,
         \R[8][21] , \R[8][20] , \R[8][19] , \R[8][18] , \R[8][17] ,
         \R[8][16] , \R[8][15] , \R[8][14] , \R[8][13] , \R[8][12] ,
         \R[8][11] , \R[8][10] , \R[8][9] , \R[8][8] , \R[8][7] , \R[8][6] ,
         \R[8][5] , \R[8][4] , \R[8][3] , \R[8][2] , \R[8][1] , \R[8][0] ,
         \R[9][31] , \R[9][30] , \R[9][29] , \R[9][28] , \R[9][27] ,
         \R[9][26] , \R[9][25] , \R[9][24] , \R[9][23] , \R[9][22] ,
         \R[9][21] , \R[9][20] , \R[9][19] , \R[9][18] , \R[9][17] ,
         \R[9][16] , \R[9][15] , \R[9][14] , \R[9][13] , \R[9][12] ,
         \R[9][11] , \R[9][10] , \R[9][9] , \R[9][8] , \R[9][7] , \R[9][6] ,
         \R[9][5] , \R[9][4] , \R[9][3] , \R[9][2] , \R[9][1] , \R[9][0] ,
         \R[10][31] , \R[10][30] , \R[10][29] , \R[10][28] , \R[10][27] ,
         \R[10][26] , \R[10][25] , \R[10][24] , \R[10][23] , \R[10][22] ,
         \R[10][21] , \R[10][20] , \R[10][19] , \R[10][18] , \R[10][17] ,
         \R[10][16] , \R[10][15] , \R[10][14] , \R[10][13] , \R[10][12] ,
         \R[10][11] , \R[10][10] , \R[10][9] , \R[10][8] , \R[10][7] ,
         \R[10][6] , \R[10][5] , \R[10][4] , \R[10][3] , \R[10][2] ,
         \R[10][1] , \R[10][0] , \R[11][31] , \R[11][30] , \R[11][29] ,
         \R[11][28] , \R[11][27] , \R[11][26] , \R[11][25] , \R[11][24] ,
         \R[11][23] , \R[11][22] , \R[11][21] , \R[11][20] , \R[11][19] ,
         \R[11][18] , \R[11][17] , \R[11][16] , \R[11][15] , \R[11][14] ,
         \R[11][13] , \R[11][12] , \R[11][11] , \R[11][10] , \R[11][9] ,
         \R[11][8] , \R[11][7] , \R[11][6] , \R[11][5] , \R[11][4] ,
         \R[11][3] , \R[11][2] , \R[11][1] , \R[11][0] , \R[12][31] ,
         \R[12][30] , \R[12][29] , \R[12][28] , \R[12][27] , \R[12][26] ,
         \R[12][25] , \R[12][24] , \R[12][23] , \R[12][22] , \R[12][21] ,
         \R[12][20] , \R[12][19] , \R[12][18] , \R[12][17] , \R[12][16] ,
         \R[12][15] , \R[12][14] , \R[12][13] , \R[12][12] , \R[12][11] ,
         \R[12][10] , \R[12][9] , \R[12][8] , \R[12][7] , \R[12][6] ,
         \R[12][5] , \R[12][4] , \R[12][3] , \R[12][2] , \R[12][1] ,
         \R[12][0] , \R[13][31] , \R[13][30] , \R[13][29] , \R[13][28] ,
         \R[13][27] , \R[13][26] , \R[13][25] , \R[13][24] , \R[13][23] ,
         \R[13][22] , \R[13][21] , \R[13][20] , \R[13][19] , \R[13][18] ,
         \R[13][17] , \R[13][16] , \R[13][15] , \R[13][14] , \R[13][13] ,
         \R[13][12] , \R[13][11] , \R[13][10] , \R[13][9] , \R[13][8] ,
         \R[13][7] , \R[13][6] , \R[13][5] , \R[13][4] , \R[13][3] ,
         \R[13][2] , \R[13][1] , \R[13][0] , \R[14][31] , \R[14][30] ,
         \R[14][29] , \R[14][28] , \R[14][27] , \R[14][26] , \R[14][25] ,
         \R[14][24] , \R[14][23] , \R[14][22] , \R[14][21] , \R[14][20] ,
         \R[14][19] , \R[14][18] , \R[14][17] , \R[14][16] , \R[14][15] ,
         \R[14][14] , \R[14][13] , \R[14][12] , \R[14][11] , \R[14][10] ,
         \R[14][9] , \R[14][8] , \R[14][7] , \R[14][6] , \R[14][5] ,
         \R[14][4] , \R[14][3] , \R[14][2] , \R[14][1] , \R[14][0] ,
         \R[15][31] , \R[15][30] , \R[15][29] , \R[15][28] , \R[15][27] ,
         \R[15][26] , \R[15][25] , \R[15][24] , \R[15][23] , \R[15][22] ,
         \R[15][21] , \R[15][20] , \R[15][19] , \R[15][18] , \R[15][17] ,
         \R[15][16] , \R[15][15] , \R[15][14] , \R[15][13] , \R[15][12] ,
         \R[15][11] , \R[15][10] , \R[15][9] , \R[15][8] , \R[15][7] ,
         \R[15][6] , \R[15][5] , \R[15][4] , \R[15][3] , \R[15][2] ,
         \R[15][1] , \R[15][0] , \R[16][31] , \R[16][30] , \R[16][29] ,
         \R[16][28] , \R[16][27] , \R[16][26] , \R[16][25] , \R[16][24] ,
         \R[16][23] , \R[16][22] , \R[16][21] , \R[16][20] , \R[16][19] ,
         \R[16][18] , \R[16][17] , \R[16][16] , \R[16][15] , \R[16][14] ,
         \R[16][13] , \R[16][12] , \R[16][11] , \R[16][10] , \R[16][9] ,
         \R[16][8] , \R[16][7] , \R[16][6] , \R[16][5] , \R[16][4] ,
         \R[16][3] , \R[16][2] , \R[16][1] , \R[16][0] , \R[17][31] ,
         \R[17][30] , \R[17][29] , \R[17][28] , \R[17][27] , \R[17][26] ,
         \R[17][25] , \R[17][24] , \R[17][23] , \R[17][22] , \R[17][21] ,
         \R[17][20] , \R[17][19] , \R[17][18] , \R[17][17] , \R[17][16] ,
         \R[17][15] , \R[17][14] , \R[17][13] , \R[17][12] , \R[17][11] ,
         \R[17][10] , \R[17][9] , \R[17][8] , \R[17][7] , \R[17][6] ,
         \R[17][5] , \R[17][4] , \R[17][3] , \R[17][2] , \R[17][1] ,
         \R[17][0] , \R[18][31] , \R[18][30] , \R[18][29] , \R[18][28] ,
         \R[18][27] , \R[18][26] , \R[18][25] , \R[18][24] , \R[18][23] ,
         \R[18][22] , \R[18][21] , \R[18][20] , \R[18][19] , \R[18][18] ,
         \R[18][17] , \R[18][16] , \R[18][15] , \R[18][14] , \R[18][13] ,
         \R[18][12] , \R[18][11] , \R[18][10] , \R[18][9] , \R[18][8] ,
         \R[18][7] , \R[18][6] , \R[18][5] , \R[18][4] , \R[18][3] ,
         \R[18][2] , \R[18][1] , \R[18][0] , \R[19][31] , \R[19][30] ,
         \R[19][29] , \R[19][28] , \R[19][27] , \R[19][26] , \R[19][25] ,
         \R[19][24] , \R[19][23] , \R[19][22] , \R[19][21] , \R[19][20] ,
         \R[19][19] , \R[19][18] , \R[19][17] , \R[19][16] , \R[19][15] ,
         \R[19][14] , \R[19][13] , \R[19][12] , \R[19][11] , \R[19][10] ,
         \R[19][9] , \R[19][8] , \R[19][7] , \R[19][6] , \R[19][5] ,
         \R[19][4] , \R[19][3] , \R[19][2] , \R[19][1] , \R[19][0] ,
         \R[20][31] , \R[20][30] , \R[20][29] , \R[20][28] , \R[20][27] ,
         \R[20][26] , \R[20][25] , \R[20][24] , \R[20][23] , \R[20][22] ,
         \R[20][21] , \R[20][20] , \R[20][19] , \R[20][18] , \R[20][17] ,
         \R[20][16] , \R[20][15] , \R[20][14] , \R[20][13] , \R[20][12] ,
         \R[20][11] , \R[20][10] , \R[20][9] , \R[20][8] , \R[20][7] ,
         \R[20][6] , \R[20][5] , \R[20][4] , \R[20][3] , \R[20][2] ,
         \R[20][1] , \R[20][0] , \R[21][31] , \R[21][30] , \R[21][29] ,
         \R[21][28] , \R[21][27] , \R[21][26] , \R[21][25] , \R[21][24] ,
         \R[21][23] , \R[21][22] , \R[21][21] , \R[21][20] , \R[21][19] ,
         \R[21][18] , \R[21][17] , \R[21][16] , \R[21][15] , \R[21][14] ,
         \R[21][13] , \R[21][12] , \R[21][11] , \R[21][10] , \R[21][9] ,
         \R[21][8] , \R[21][7] , \R[21][6] , \R[21][5] , \R[21][4] ,
         \R[21][3] , \R[21][2] , \R[21][1] , \R[21][0] , \R[22][31] ,
         \R[22][30] , \R[22][29] , \R[22][28] , \R[22][27] , \R[22][26] ,
         \R[22][25] , \R[22][24] , \R[22][23] , \R[22][22] , \R[22][21] ,
         \R[22][20] , \R[22][19] , \R[22][18] , \R[22][17] , \R[22][16] ,
         \R[22][15] , \R[22][14] , \R[22][13] , \R[22][12] , \R[22][11] ,
         \R[22][10] , \R[22][9] , \R[22][8] , \R[22][7] , \R[22][6] ,
         \R[22][5] , \R[22][4] , \R[22][3] , \R[22][2] , \R[22][1] ,
         \R[22][0] , \R[23][31] , \R[23][30] , \R[23][29] , \R[23][28] ,
         \R[23][27] , \R[23][26] , \R[23][25] , \R[23][24] , \R[23][23] ,
         \R[23][22] , \R[23][21] , \R[23][20] , \R[23][19] , \R[23][18] ,
         \R[23][17] , \R[23][16] , \R[23][15] , \R[23][14] , \R[23][13] ,
         \R[23][12] , \R[23][11] , \R[23][10] , \R[23][9] , \R[23][8] ,
         \R[23][7] , \R[23][6] , \R[23][5] , \R[23][4] , \R[23][3] ,
         \R[23][2] , \R[23][1] , \R[23][0] , \R[24][31] , \R[24][30] ,
         \R[24][29] , \R[24][28] , \R[24][27] , \R[24][26] , \R[24][25] ,
         \R[24][24] , \R[24][23] , \R[24][22] , \R[24][21] , \R[24][20] ,
         \R[24][19] , \R[24][18] , \R[24][17] , \R[24][16] , \R[24][15] ,
         \R[24][14] , \R[24][13] , \R[24][12] , \R[24][11] , \R[24][10] ,
         \R[24][9] , \R[24][8] , \R[24][7] , \R[24][6] , \R[24][5] ,
         \R[24][4] , \R[24][3] , \R[24][2] , \R[24][1] , \R[24][0] ,
         \R[25][31] , \R[25][30] , \R[25][29] , \R[25][28] , \R[25][27] ,
         \R[25][26] , \R[25][25] , \R[25][24] , \R[25][23] , \R[25][22] ,
         \R[25][21] , \R[25][20] , \R[25][19] , \R[25][18] , \R[25][17] ,
         \R[25][16] , \R[25][15] , \R[25][14] , \R[25][13] , \R[25][12] ,
         \R[25][11] , \R[25][10] , \R[25][9] , \R[25][8] , \R[25][7] ,
         \R[25][6] , \R[25][5] , \R[25][4] , \R[25][3] , \R[25][2] ,
         \R[25][1] , \R[25][0] , \R[26][31] , \R[26][30] , \R[26][29] ,
         \R[26][28] , \R[26][27] , \R[26][26] , \R[26][25] , \R[26][24] ,
         \R[26][23] , \R[26][22] , \R[26][21] , \R[26][20] , \R[26][19] ,
         \R[26][18] , \R[26][17] , \R[26][16] , \R[26][15] , \R[26][14] ,
         \R[26][13] , \R[26][12] , \R[26][11] , \R[26][10] , \R[26][9] ,
         \R[26][8] , \R[26][7] , \R[26][6] , \R[26][5] , \R[26][4] ,
         \R[26][3] , \R[26][2] , \R[26][1] , \R[26][0] , \R[27][31] ,
         \R[27][30] , \R[27][29] , \R[27][28] , \R[27][27] , \R[27][26] ,
         \R[27][25] , \R[27][24] , \R[27][23] , \R[27][22] , \R[27][21] ,
         \R[27][20] , \R[27][19] , \R[27][18] , \R[27][17] , \R[27][16] ,
         \R[27][15] , \R[27][14] , \R[27][13] , \R[27][12] , \R[27][11] ,
         \R[27][10] , \R[27][9] , \R[27][8] , \R[27][7] , \R[27][6] ,
         \R[27][5] , \R[27][4] , \R[27][3] , \R[27][2] , \R[27][1] ,
         \R[27][0] , \R[28][31] , \R[28][30] , \R[28][29] , \R[28][28] ,
         \R[28][27] , \R[28][26] , \R[28][25] , \R[28][24] , \R[28][23] ,
         \R[28][22] , \R[28][21] , \R[28][20] , \R[28][19] , \R[28][18] ,
         \R[28][17] , \R[28][16] , \R[28][15] , \R[28][14] , \R[28][13] ,
         \R[28][12] , \R[28][11] , \R[28][10] , \R[28][9] , \R[28][8] ,
         \R[28][7] , \R[28][6] , \R[28][5] , \R[28][4] , \R[28][3] ,
         \R[28][2] , \R[28][1] , \R[28][0] , \R[29][31] , \R[29][30] ,
         \R[29][29] , \R[29][28] , \R[29][27] , \R[29][26] , \R[29][25] ,
         \R[29][24] , \R[29][23] , \R[29][22] , \R[29][21] , \R[29][20] ,
         \R[29][19] , \R[29][18] , \R[29][17] , \R[29][16] , \R[29][15] ,
         \R[29][14] , \R[29][13] , \R[29][12] , \R[29][11] , \R[29][10] ,
         \R[29][9] , \R[29][8] , \R[29][7] , \R[29][6] , \R[29][5] ,
         \R[29][4] , \R[29][3] , \R[29][2] , \R[29][1] , \R[29][0] ,
         \R[30][31] , \R[30][30] , \R[30][29] , \R[30][28] , \R[30][27] ,
         \R[30][26] , \R[30][25] , \R[30][24] , \R[30][23] , \R[30][22] ,
         \R[30][21] , \R[30][20] , \R[30][19] , \R[30][18] , \R[30][17] ,
         \R[30][16] , \R[30][15] , \R[30][14] , \R[30][13] , \R[30][12] ,
         \R[30][11] , \R[30][10] , \R[30][9] , \R[30][8] , \R[30][7] ,
         \R[30][6] , \R[30][5] , \R[30][4] , \R[30][3] , \R[30][2] ,
         \R[30][1] , \R[30][0] , \R[31][31] , \R[31][30] , \R[31][29] ,
         \R[31][28] , \R[31][27] , \R[31][26] , \R[31][25] , \R[31][24] ,
         \R[31][23] , \R[31][22] , \R[31][21] , \R[31][20] , \R[31][19] ,
         \R[31][18] , \R[31][17] , \R[31][16] , \R[31][15] , \R[31][14] ,
         \R[31][13] , \R[31][12] , \R[31][11] , \R[31][10] , \R[31][9] ,
         \R[31][8] , \R[31][7] , \R[31][6] , \R[31][5] , \R[31][4] ,
         \R[31][3] , \R[31][2] , \R[31][1] , \R[31][0] , N60, N61, N62, N63,
         N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77,
         N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91,
         N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, N136,
         N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147,
         N148, N149, N150, N151, N152, N153, N154, N155, N156, N157,
         \seIM[31] , N190, N192, N193, N195, N197, N198, N199, N200, N203,
         N204, N205, N207, N208, N217, N218, N219, N220, N222, N223, N224,
         N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235,
         N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, N246,
         N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N257,
         N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268,
         N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, N279,
         N280, N281, N282, N283, N284, N285, N401, N402, N403, N404, N405,
         N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416,
         N417, N418, N419, N420, N421, N422, N423, N424, N425, N426, N427,
         N428, N429, N430, N431, N432, N433, N434, N435, N436, N437, N438,
         N439, N440, N441, N442, N443, N444, N445, N446, N447, N448, N449,
         N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460,
         N461, N462, N463, N464, N593, N594, N595, N596, N597, N598, N599,
         N600, N601, N602, N603, N604, N605, N606, N607, N608, N609, N610,
         N611, N612, N613, N614, N615, N616, N617, N618, N619, N620, N621,
         N622, N623, N624, N657, N658, N659, N660, N661, N662, N663, N664,
         N665, N666, N667, N668, N669, N670, N671, N672, N673, N674, N675,
         N676, N677, N678, N679, N680, N681, N682, N683, N684, N685, N686,
         N687, N688, N785, N786, N787, N788, N789, N790, N791, N792, N793,
         N794, N795, N796, N797, N798, N799, N800, N801, N802, N803, N804,
         N805, N806, N807, N808, N809, N810, N811, N812, N813, N814, N815,
         N816, N864, N865, N866, N867, N868, N869, N870, N871, N872, N873,
         N874, N875, N876, N877, N878, N879, N880, N881, N882, N883, N884,
         N885, N886, N887, N888, N889, N890, N891, N892, N893, N894, N895,
         N896, N897, N898, N899, N900, N901, N902, N903, N904, N905, N906,
         N907, N908, N909, N910, N911, N912, N913, N914, N915, N916, N917,
         N918, N919, N920, N921, N922, N923, N924, N925, N926, N927, N928,
         N929, N930, N931, N932, N933, N934, N935, N936, N937, N938, N939,
         N940, N941, N942, N943, N944, N945, N946, N947, N948, N949, N950,
         N951, N952, N953, N954, N955, N956, N957, N958, N959, N960, N993,
         N994, N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003, N1004,
         N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013, N1014,
         N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023, N1024,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n78, n111, n113, n114,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n151, n152, n154, n155, n156, n158, n159, n161, n163, n164,
         n165, n167, n168, n170, n171, n173, n175, n177, n179, n180, n181,
         n183, n184, n186, n188, n190, n191, n193, n194, n196, n198, n201,
         n203, n204, n206, n207, n209, n211, n213, n214, n216, n217, n219,
         n222, n225, n228, n229, n230, n231, n232, n233, n234, n235, n237,
         n238, n239, n240, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n518, n519, n520, n521, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n543, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646,
         N645, N644, N643, N642,
         \sub_1_root_add_0_root_add_137_ni_b0/carry[2] ,
         \sub_1_root_add_0_root_add_137_ni_b0/carry[3] ,
         \sub_1_root_add_0_root_add_137_ni_b0/carry[4] ,
         \sub_1_root_add_0_root_add_137_ni_b0/carry[5] ,
         \sub_1_root_add_0_root_add_137_ni_b0/carry[6] ,
         \sub_1_root_add_0_root_add_137_ni_b0/carry[7] ,
         \sub_1_root_add_0_root_add_137_ni_b0/carry[8] ,
         \sub_1_root_add_0_root_add_137_ni_b0/carry[9] ,
         \sub_1_root_add_0_root_add_137_ni_b0/carry[10] ,
         \sub_1_root_add_0_root_add_137_ni_b0/carry[11] ,
         \sub_1_root_add_0_root_add_137_ni_b0/carry[12] ,
         \sub_1_root_add_0_root_add_137_ni_b0/carry[13] ,
         \sub_1_root_add_0_root_add_137_ni_b0/carry[14] , n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045;
  wire   [31:0] counter;
  assign N46 = instruction[15];
  assign N47 = instruction[16];
  assign N48 = instruction[17];
  assign N49 = instruction[18];
  assign N50 = instruction[19];
  assign N51 = instruction[10];
  assign N52 = instruction[11];
  assign N53 = instruction[12];
  assign N54 = instruction[13];
  assign \seIM[31]  = instruction[14];
  assign N656 = instruction[0];

  SingleCycleProcessor_DW_cmp_0 lt_182 ( .A({N190, n2652, N192, N193, n2651, 
        N195, n2650, N197, N198, N199, N200, n2648, n2649, N203, N204, N205, 
        n2653, N207, N208, n2677, n2676, n2673, n2674, n2675, n2671, n2672, 
        n2655, N217, N218, N219, N220, n2670}), .B({N222, N223, N224, N225, 
        N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, 
        N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, 
        N250, N251, N252, N253}), .TC(1'b1), .GE_LT(1'b1), .GE_GT_EQ(1'b0), 
        .GE_LT_GT_LE(N960) );
  SingleCycleProcessor_DW_leftsh_0 sll_169 ( .A({N190, n2652, N192, N193, 
        n2651, N195, n2650, N197, N198, N199, N200, n2648, n2649, N203, N204, 
        N205, n2653, N207, N208, n2677, n2676, n2673, n2674, n2675, n2671, 
        n2672, n2655, N217, N218, N219, N220, n2670}), .SH({instruction[4:1], 
        N656}), .B({N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, 
        N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, 
        N937, N936, N935, N934, N933, N932, N931, N930, N929, N928}) );
  SingleCycleProcessor_DW_rightsh_0 srl_165 ( .A({N190, n2652, N192, N193, 
        n2651, N195, n2650, N197, N198, N199, N200, n2648, n2649, N203, N204, 
        N205, n2653, N207, N208, n2677, n2676, n2673, n2674, n2675, n2671, 
        n2672, n2655, N217, N218, N219, N220, n2670}), .DATA_TC(1'b0), .SH({
        instruction[4:1], N656}), .B({N927, N926, N925, N924, N923, N922, N921, 
        N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, 
        N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, 
        N896}) );
  SingleCycleProcessor_DW01_add_0 add_1_root_add_157_2 ( .A({N190, n2652, N192, 
        N193, n2651, N195, n2650, N197, N198, N199, N200, n2648, n2649, N203, 
        N204, N205, n2653, N207, N208, n2677, n2676, n2673, n2674, n2675, 
        n2671, n2672, n2655, N217, N218, N219, N220, n2670}), .B({1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, n3972, n3978, n3979, n3981, n3982, n4040, n4041, 
        n4042, n4043, n4044, n3977, n3976, n3975, n3974, n3787}), .CI(1'b1), 
        .SUM({N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, 
        N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, 
        N872, N871, N870, N869, N868, N867, N866, N865, N864}) );
  SingleCycleProcessor_DW01_add_1 add_153 ( .A({N190, n2652, N192, N193, n2651, 
        N195, n2650, N197, N198, N199, N200, n2648, n2649, N203, N204, N205, 
        n2653, N207, N208, n2677, n2676, n2673, n2674, n2675, n2671, n2672, 
        n2655, N217, N218, N219, N220, n2670}), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, n3770, N54, N53, n3980, N51, instruction[9:1], N656}), .CI(1'b0), 
        .SUM({N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, 
        N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, 
        N793, N792, N791, N790, N789, N788, N787, N786, N785}) );
  SingleCycleProcessor_DW01_add_2 add_133 ( .A({N190, n2652, N192, N193, n2651, 
        N195, n2650, N197, N198, N199, N200, n2648, n2649, N203, N204, N205, 
        n2653, N207, N208, n2677, n2676, n2673, n2674, n2675, n2671, n2672, 
        n2655, N217, N218, N219, N220, n2663}), .B({n3770, n3770, n3770, n3767, 
        n3770, \seIM[31] , n3770, \seIM[31] , \seIM[31] , n3770, n3767, 
        \seIM[31] , n3770, \seIM[31] , n3770, \seIM[31] , n3767, n3770, N54, 
        N53, n3980, N51, instruction[9:1], N656}), .CI(1'b0), .SUM({N624, N623, 
        N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, 
        N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, 
        N598, N597, N596, N595, N594, N593}) );
  SingleCycleProcessor_DW01_sub_0 sub_113 ( .A({N190, n2652, N192, N193, n2651, 
        N195, n2650, N197, N198, N199, N200, n2648, n2649, N203, N204, N205, 
        n2653, N207, N208, n2677, n2676, n2673, n2674, n2675, n2671, n2672, 
        n2655, N217, N218, N219, N220, n2670}), .B({N222, N223, N224, N225, 
        N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, 
        N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, 
        N250, N251, N252, N253}), .CI(1'b0), .DIFF({N464, N463, N462, N461, 
        N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, 
        N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, 
        N436, N435, N434, N433}) );
  SingleCycleProcessor_DW01_add_3 add_109 ( .A({N190, n2652, N192, N193, n2651, 
        N195, n2650, N197, N198, N199, N200, n2648, n2649, N203, N204, N205, 
        n2653, N207, N208, n2677, n2676, n2673, n2674, n2675, n2671, n2672, 
        n2655, N217, N218, N219, N220, n2670}), .B({N222, N223, N224, N225, 
        N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, 
        N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, 
        N250, N251, N252, N253}), .CI(1'b0), .SUM({N432, N431, N430, N429, 
        N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, 
        N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, 
        N404, N403, N402, N401}) );
  SingleCycleProcessor_DW01_inc_0 add_57 ( .A(counter), .SUM({N91, N90, N89, 
        N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, 
        N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, 
        N60}) );
  SingleCycleProcessor_DW01_add_4 r408 ( .A(PC), .B({n3767, \seIM[31] , 
        \seIM[31] , \seIM[31] , \seIM[31] , \seIM[31] , \seIM[31] , \seIM[31] , 
        \seIM[31] , \seIM[31] , \seIM[31] , \seIM[31] , \seIM[31] , \seIM[31] , 
        \seIM[31] , \seIM[31] , \seIM[31] , \seIM[31] , N54, N53, n3980, N51, 
        instruction[9:1], N656}), .CI(1'b1), .SUM({N1024, N1023, N1022, N1021, 
        N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, 
        N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, 
        N1000, N999, N998, N997, N996, N995, N994, N993}) );
  SingleCycleProcessor_DW01_inc_1 r398 ( .A(PC), .SUM({N285, N284, N283, N282, 
        N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, 
        N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, 
        N257, N256, N255, N254}) );
  SingleCycleProcessor_DW01_add_5 add_0_root_add_0_root_add_137_ni_b0 ( .A({
        n2657, n2657, n2657, n2657, n2657, n2657, n2657, n2657, n2657, n2657, 
        n2657, n2657, n2657, n2657, n2657, n2657, n2657, N642, N643, N644, 
        N645, N646, N647, N648, N649, N650, N651, N652, N653, N654, N655, N656}), .B({N190, n2652, N192, N193, n2651, N195, n2650, N197, N198, N199, N200, 
        n2648, n2649, N203, N204, N205, n2653, N207, N208, n2677, n2676, n2673, 
        n2674, n2675, n2671, n2672, n2655, N217, N218, N219, N220, n2670}), 
        .CI(1'b0), .SUM({N688, N687, N686, N685, N684, N683, N682, N681, N680, 
        N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, 
        N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657}) );
  DFFRX1 \PC_reg[31]  ( .D(n2631), .CK(clk), .RN(reset_n), .Q(PC[31]), .QN(
        n1607) );
  DFFRX1 \PC_reg[30]  ( .D(n2630), .CK(clk), .RN(reset_n), .Q(PC[30]), .QN(
        n1596) );
  DFFRX1 \PC_reg[28]  ( .D(n2601), .CK(clk), .RN(reset_n), .Q(PC[28]), .QN(
        n1567) );
  DFFRX1 \PC_reg[29]  ( .D(n2600), .CK(clk), .RN(reset_n), .Q(PC[29]), .QN(
        n1566) );
  DFFRX1 \counter_reg[31]  ( .D(N157), .CK(clk), .RN(reset_n), .Q(counter[31]), 
        .QN(n40) );
  DFFRX1 \counter_reg[28]  ( .D(N154), .CK(clk), .RN(reset_n), .Q(counter[28]), 
        .QN(n43) );
  DFFRX1 \counter_reg[24]  ( .D(N150), .CK(clk), .RN(reset_n), .Q(counter[24]), 
        .QN(n47) );
  DFFRX1 \counter_reg[20]  ( .D(N146), .CK(clk), .RN(reset_n), .Q(counter[20]), 
        .QN(n1599) );
  DFFRX1 \counter_reg[16]  ( .D(N142), .CK(clk), .RN(reset_n), .Q(counter[16]), 
        .QN(n1603) );
  DFFRX1 \counter_reg[26]  ( .D(N152), .CK(clk), .RN(reset_n), .Q(counter[26]), 
        .QN(n45) );
  DFFRX1 \counter_reg[22]  ( .D(N148), .CK(clk), .RN(reset_n), .Q(counter[22]), 
        .QN(n1601) );
  DFFRX1 \counter_reg[18]  ( .D(N144), .CK(clk), .RN(reset_n), .Q(counter[18]), 
        .QN(n1605) );
  DFFRX1 \counter_reg[29]  ( .D(N155), .CK(clk), .RN(reset_n), .Q(counter[29]), 
        .QN(n42) );
  DFFRX1 \counter_reg[25]  ( .D(N151), .CK(clk), .RN(reset_n), .Q(counter[25]), 
        .QN(n46) );
  DFFRX1 \counter_reg[21]  ( .D(N147), .CK(clk), .RN(reset_n), .Q(counter[21]), 
        .QN(n1600) );
  DFFRX1 \counter_reg[17]  ( .D(N143), .CK(clk), .RN(reset_n), .Q(counter[17]), 
        .QN(n1604) );
  DFFRX1 \counter_reg[30]  ( .D(N156), .CK(clk), .RN(reset_n), .Q(counter[30]), 
        .QN(n41) );
  DFFRX1 \counter_reg[27]  ( .D(N153), .CK(clk), .RN(reset_n), .Q(counter[27]), 
        .QN(n44) );
  DFFRX1 \counter_reg[23]  ( .D(N149), .CK(clk), .RN(reset_n), .Q(counter[23]), 
        .QN(n1602) );
  DFFRX1 \counter_reg[19]  ( .D(N145), .CK(clk), .RN(reset_n), .Q(counter[19]), 
        .QN(n1606) );
  DFFRX1 \PC_reg[22]  ( .D(n2607), .CK(clk), .RN(reset_n), .Q(PC[22]), .QN(
        n1573) );
  DFFRX1 \PC_reg[23]  ( .D(n2606), .CK(clk), .RN(reset_n), .Q(PC[23]), .QN(
        n1572) );
  DFFRX1 \PC_reg[24]  ( .D(n2605), .CK(clk), .RN(reset_n), .Q(PC[24]), .QN(
        n1571) );
  DFFRX1 \PC_reg[25]  ( .D(n2604), .CK(clk), .RN(reset_n), .Q(PC[25]), .QN(
        n1570) );
  DFFRX1 \PC_reg[26]  ( .D(n2603), .CK(clk), .RN(reset_n), .Q(PC[26]), .QN(
        n1569) );
  DFFRX1 \PC_reg[27]  ( .D(n2602), .CK(clk), .RN(reset_n), .Q(PC[27]), .QN(
        n1568) );
  DFFRX1 \R_reg[7][24]  ( .D(n2383), .CK(clk), .RN(reset_n), .Q(\R[7][24] ), 
        .QN(n1349) );
  DFFRX1 \R_reg[7][25]  ( .D(n2382), .CK(clk), .RN(reset_n), .Q(\R[7][25] ), 
        .QN(n1348) );
  DFFRX1 \R_reg[7][26]  ( .D(n2381), .CK(clk), .RN(reset_n), .Q(\R[7][26] ), 
        .QN(n1347) );
  DFFRX1 \R_reg[7][27]  ( .D(n2380), .CK(clk), .RN(reset_n), .Q(\R[7][27] ), 
        .QN(n1346) );
  DFFRX1 \R_reg[7][28]  ( .D(n2379), .CK(clk), .RN(reset_n), .Q(\R[7][28] ), 
        .QN(n1345) );
  DFFRX1 \R_reg[7][29]  ( .D(n2378), .CK(clk), .RN(reset_n), .Q(\R[7][29] ), 
        .QN(n1344) );
  DFFRX1 \R_reg[7][30]  ( .D(n2377), .CK(clk), .RN(reset_n), .Q(\R[7][30] ), 
        .QN(n1343) );
  DFFRX1 \R_reg[7][31]  ( .D(n2376), .CK(clk), .RN(reset_n), .Q(\R[7][31] ), 
        .QN(n1342) );
  DFFRX1 \R_reg[11][24]  ( .D(n2255), .CK(clk), .RN(reset_n), .Q(\R[11][24] ), 
        .QN(n1221) );
  DFFRX1 \R_reg[11][25]  ( .D(n2254), .CK(clk), .RN(reset_n), .Q(\R[11][25] ), 
        .QN(n1220) );
  DFFRX1 \R_reg[11][26]  ( .D(n2253), .CK(clk), .RN(reset_n), .Q(\R[11][26] ), 
        .QN(n1219) );
  DFFRX1 \R_reg[11][27]  ( .D(n2252), .CK(clk), .RN(reset_n), .Q(\R[11][27] ), 
        .QN(n1218) );
  DFFRX1 \R_reg[11][28]  ( .D(n2251), .CK(clk), .RN(reset_n), .Q(\R[11][28] ), 
        .QN(n1217) );
  DFFRX1 \R_reg[11][29]  ( .D(n2250), .CK(clk), .RN(reset_n), .Q(\R[11][29] ), 
        .QN(n1216) );
  DFFRX1 \R_reg[11][30]  ( .D(n2249), .CK(clk), .RN(reset_n), .Q(\R[11][30] ), 
        .QN(n1215) );
  DFFRX1 \R_reg[11][31]  ( .D(n2248), .CK(clk), .RN(reset_n), .Q(\R[11][31] ), 
        .QN(n1214) );
  DFFRX1 \R_reg[15][24]  ( .D(n2127), .CK(clk), .RN(reset_n), .Q(\R[15][24] ), 
        .QN(n1093) );
  DFFRX1 \R_reg[15][25]  ( .D(n2126), .CK(clk), .RN(reset_n), .Q(\R[15][25] ), 
        .QN(n1092) );
  DFFRX1 \R_reg[15][26]  ( .D(n2125), .CK(clk), .RN(reset_n), .Q(\R[15][26] ), 
        .QN(n1091) );
  DFFRX1 \R_reg[15][27]  ( .D(n2124), .CK(clk), .RN(reset_n), .Q(\R[15][27] ), 
        .QN(n1090) );
  DFFRX1 \R_reg[15][28]  ( .D(n2123), .CK(clk), .RN(reset_n), .Q(\R[15][28] ), 
        .QN(n1089) );
  DFFRX1 \R_reg[15][29]  ( .D(n2122), .CK(clk), .RN(reset_n), .Q(\R[15][29] ), 
        .QN(n1088) );
  DFFRX1 \R_reg[15][30]  ( .D(n2121), .CK(clk), .RN(reset_n), .Q(\R[15][30] ), 
        .QN(n1087) );
  DFFRX1 \R_reg[15][31]  ( .D(n2120), .CK(clk), .RN(reset_n), .Q(\R[15][31] ), 
        .QN(n1086) );
  DFFRX1 \R_reg[19][24]  ( .D(n1999), .CK(clk), .RN(reset_n), .Q(\R[19][24] ), 
        .QN(n965) );
  DFFRX1 \R_reg[19][25]  ( .D(n1998), .CK(clk), .RN(reset_n), .Q(\R[19][25] ), 
        .QN(n964) );
  DFFRX1 \R_reg[19][26]  ( .D(n1997), .CK(clk), .RN(reset_n), .Q(\R[19][26] ), 
        .QN(n963) );
  DFFRX1 \R_reg[19][27]  ( .D(n1996), .CK(clk), .RN(reset_n), .Q(\R[19][27] ), 
        .QN(n962) );
  DFFRX1 \R_reg[19][28]  ( .D(n1995), .CK(clk), .RN(reset_n), .Q(\R[19][28] ), 
        .QN(n961) );
  DFFRX1 \R_reg[19][29]  ( .D(n1994), .CK(clk), .RN(reset_n), .Q(\R[19][29] ), 
        .QN(n960) );
  DFFRX1 \R_reg[19][30]  ( .D(n1993), .CK(clk), .RN(reset_n), .Q(\R[19][30] ), 
        .QN(n959) );
  DFFRX1 \R_reg[19][31]  ( .D(n1992), .CK(clk), .RN(reset_n), .Q(\R[19][31] ), 
        .QN(n958) );
  DFFRX1 \R_reg[23][24]  ( .D(n1871), .CK(clk), .RN(reset_n), .Q(\R[23][24] ), 
        .QN(n837) );
  DFFRX1 \R_reg[23][25]  ( .D(n1870), .CK(clk), .RN(reset_n), .Q(\R[23][25] ), 
        .QN(n836) );
  DFFRX1 \R_reg[23][26]  ( .D(n1869), .CK(clk), .RN(reset_n), .Q(\R[23][26] ), 
        .QN(n835) );
  DFFRX1 \R_reg[23][27]  ( .D(n1868), .CK(clk), .RN(reset_n), .Q(\R[23][27] ), 
        .QN(n834) );
  DFFRX1 \R_reg[23][28]  ( .D(n1867), .CK(clk), .RN(reset_n), .Q(\R[23][28] ), 
        .QN(n833) );
  DFFRX1 \R_reg[23][29]  ( .D(n1866), .CK(clk), .RN(reset_n), .Q(\R[23][29] ), 
        .QN(n832) );
  DFFRX1 \R_reg[23][30]  ( .D(n1865), .CK(clk), .RN(reset_n), .Q(\R[23][30] ), 
        .QN(n831) );
  DFFRX1 \R_reg[23][31]  ( .D(n1864), .CK(clk), .RN(reset_n), .Q(\R[23][31] ), 
        .QN(n830) );
  DFFRX1 \R_reg[27][24]  ( .D(n1743), .CK(clk), .RN(reset_n), .Q(\R[27][24] ), 
        .QN(n709) );
  DFFRX1 \R_reg[27][25]  ( .D(n1742), .CK(clk), .RN(reset_n), .Q(\R[27][25] ), 
        .QN(n708) );
  DFFRX1 \R_reg[27][26]  ( .D(n1741), .CK(clk), .RN(reset_n), .Q(\R[27][26] ), 
        .QN(n707) );
  DFFRX1 \R_reg[27][27]  ( .D(n1740), .CK(clk), .RN(reset_n), .Q(\R[27][27] ), 
        .QN(n706) );
  DFFRX1 \R_reg[27][28]  ( .D(n1739), .CK(clk), .RN(reset_n), .Q(\R[27][28] ), 
        .QN(n705) );
  DFFRX1 \R_reg[27][29]  ( .D(n1738), .CK(clk), .RN(reset_n), .Q(\R[27][29] ), 
        .QN(n704) );
  DFFRX1 \R_reg[27][30]  ( .D(n1737), .CK(clk), .RN(reset_n), .Q(\R[27][30] ), 
        .QN(n703) );
  DFFRX1 \R_reg[27][31]  ( .D(n1736), .CK(clk), .RN(reset_n), .Q(\R[27][31] ), 
        .QN(n702) );
  DFFRX1 \R_reg[31][24]  ( .D(n1615), .CK(clk), .RN(reset_n), .Q(\R[31][24] ), 
        .QN(n581) );
  DFFRX1 \R_reg[31][25]  ( .D(n1614), .CK(clk), .RN(reset_n), .Q(\R[31][25] ), 
        .QN(n580) );
  DFFRX1 \R_reg[31][26]  ( .D(n1613), .CK(clk), .RN(reset_n), .Q(\R[31][26] ), 
        .QN(n579) );
  DFFRX1 \R_reg[31][27]  ( .D(n1612), .CK(clk), .RN(reset_n), .Q(\R[31][27] ), 
        .QN(n578) );
  DFFRX1 \R_reg[31][28]  ( .D(n1611), .CK(clk), .RN(reset_n), .Q(\R[31][28] ), 
        .QN(n577) );
  DFFRX1 \R_reg[31][29]  ( .D(n1610), .CK(clk), .RN(reset_n), .Q(\R[31][29] ), 
        .QN(n576) );
  DFFRX1 \R_reg[31][30]  ( .D(n1609), .CK(clk), .RN(reset_n), .Q(\R[31][30] ), 
        .QN(n575) );
  DFFRX1 \R_reg[31][31]  ( .D(n1608), .CK(clk), .RN(reset_n), .Q(\R[31][31] ), 
        .QN(n574) );
  DFFRX1 \R_reg[5][24]  ( .D(n2447), .CK(clk), .RN(reset_n), .Q(\R[5][24] ), 
        .QN(n1413) );
  DFFRX1 \R_reg[5][25]  ( .D(n2446), .CK(clk), .RN(reset_n), .Q(\R[5][25] ), 
        .QN(n1412) );
  DFFRX1 \R_reg[5][26]  ( .D(n2445), .CK(clk), .RN(reset_n), .Q(\R[5][26] ), 
        .QN(n1411) );
  DFFRX1 \R_reg[5][27]  ( .D(n2444), .CK(clk), .RN(reset_n), .Q(\R[5][27] ), 
        .QN(n1410) );
  DFFRX1 \R_reg[5][28]  ( .D(n2443), .CK(clk), .RN(reset_n), .Q(\R[5][28] ), 
        .QN(n1409) );
  DFFRX1 \R_reg[5][29]  ( .D(n2442), .CK(clk), .RN(reset_n), .Q(\R[5][29] ), 
        .QN(n1408) );
  DFFRX1 \R_reg[5][30]  ( .D(n2441), .CK(clk), .RN(reset_n), .Q(\R[5][30] ), 
        .QN(n1407) );
  DFFRX1 \R_reg[5][31]  ( .D(n2440), .CK(clk), .RN(reset_n), .Q(\R[5][31] ), 
        .QN(n1406) );
  DFFRX1 \R_reg[9][24]  ( .D(n2319), .CK(clk), .RN(reset_n), .Q(\R[9][24] ), 
        .QN(n1285) );
  DFFRX1 \R_reg[9][25]  ( .D(n2318), .CK(clk), .RN(reset_n), .Q(\R[9][25] ), 
        .QN(n1284) );
  DFFRX1 \R_reg[9][26]  ( .D(n2317), .CK(clk), .RN(reset_n), .Q(\R[9][26] ), 
        .QN(n1283) );
  DFFRX1 \R_reg[9][27]  ( .D(n2316), .CK(clk), .RN(reset_n), .Q(\R[9][27] ), 
        .QN(n1282) );
  DFFRX1 \R_reg[9][28]  ( .D(n2315), .CK(clk), .RN(reset_n), .Q(\R[9][28] ), 
        .QN(n1281) );
  DFFRX1 \R_reg[9][29]  ( .D(n2314), .CK(clk), .RN(reset_n), .Q(\R[9][29] ), 
        .QN(n1280) );
  DFFRX1 \R_reg[9][30]  ( .D(n2313), .CK(clk), .RN(reset_n), .Q(\R[9][30] ), 
        .QN(n1279) );
  DFFRX1 \R_reg[9][31]  ( .D(n2312), .CK(clk), .RN(reset_n), .Q(\R[9][31] ), 
        .QN(n1278) );
  DFFRX1 \R_reg[13][24]  ( .D(n2191), .CK(clk), .RN(reset_n), .Q(\R[13][24] ), 
        .QN(n1157) );
  DFFRX1 \R_reg[13][25]  ( .D(n2190), .CK(clk), .RN(reset_n), .Q(\R[13][25] ), 
        .QN(n1156) );
  DFFRX1 \R_reg[13][26]  ( .D(n2189), .CK(clk), .RN(reset_n), .Q(\R[13][26] ), 
        .QN(n1155) );
  DFFRX1 \R_reg[13][27]  ( .D(n2188), .CK(clk), .RN(reset_n), .Q(\R[13][27] ), 
        .QN(n1154) );
  DFFRX1 \R_reg[13][28]  ( .D(n2187), .CK(clk), .RN(reset_n), .Q(\R[13][28] ), 
        .QN(n1153) );
  DFFRX1 \R_reg[13][29]  ( .D(n2186), .CK(clk), .RN(reset_n), .Q(\R[13][29] ), 
        .QN(n1152) );
  DFFRX1 \R_reg[13][30]  ( .D(n2185), .CK(clk), .RN(reset_n), .Q(\R[13][30] ), 
        .QN(n1151) );
  DFFRX1 \R_reg[13][31]  ( .D(n2184), .CK(clk), .RN(reset_n), .Q(\R[13][31] ), 
        .QN(n1150) );
  DFFRX1 \R_reg[17][24]  ( .D(n2063), .CK(clk), .RN(reset_n), .Q(\R[17][24] ), 
        .QN(n1029) );
  DFFRX1 \R_reg[17][25]  ( .D(n2062), .CK(clk), .RN(reset_n), .Q(\R[17][25] ), 
        .QN(n1028) );
  DFFRX1 \R_reg[17][26]  ( .D(n2061), .CK(clk), .RN(reset_n), .Q(\R[17][26] ), 
        .QN(n1027) );
  DFFRX1 \R_reg[17][27]  ( .D(n2060), .CK(clk), .RN(reset_n), .Q(\R[17][27] ), 
        .QN(n1026) );
  DFFRX1 \R_reg[17][28]  ( .D(n2059), .CK(clk), .RN(reset_n), .Q(\R[17][28] ), 
        .QN(n1025) );
  DFFRX1 \R_reg[17][29]  ( .D(n2058), .CK(clk), .RN(reset_n), .Q(\R[17][29] ), 
        .QN(n1024) );
  DFFRX1 \R_reg[17][30]  ( .D(n2057), .CK(clk), .RN(reset_n), .Q(\R[17][30] ), 
        .QN(n1023) );
  DFFRX1 \R_reg[17][31]  ( .D(n2056), .CK(clk), .RN(reset_n), .Q(\R[17][31] ), 
        .QN(n1022) );
  DFFRX1 \R_reg[21][24]  ( .D(n1935), .CK(clk), .RN(reset_n), .Q(\R[21][24] ), 
        .QN(n901) );
  DFFRX1 \R_reg[21][25]  ( .D(n1934), .CK(clk), .RN(reset_n), .Q(\R[21][25] ), 
        .QN(n900) );
  DFFRX1 \R_reg[21][26]  ( .D(n1933), .CK(clk), .RN(reset_n), .Q(\R[21][26] ), 
        .QN(n899) );
  DFFRX1 \R_reg[21][27]  ( .D(n1932), .CK(clk), .RN(reset_n), .Q(\R[21][27] ), 
        .QN(n898) );
  DFFRX1 \R_reg[21][28]  ( .D(n1931), .CK(clk), .RN(reset_n), .Q(\R[21][28] ), 
        .QN(n897) );
  DFFRX1 \R_reg[21][29]  ( .D(n1930), .CK(clk), .RN(reset_n), .Q(\R[21][29] ), 
        .QN(n896) );
  DFFRX1 \R_reg[21][30]  ( .D(n1929), .CK(clk), .RN(reset_n), .Q(\R[21][30] ), 
        .QN(n895) );
  DFFRX1 \R_reg[21][31]  ( .D(n1928), .CK(clk), .RN(reset_n), .Q(\R[21][31] ), 
        .QN(n894) );
  DFFRX1 \R_reg[25][24]  ( .D(n1807), .CK(clk), .RN(reset_n), .Q(\R[25][24] ), 
        .QN(n773) );
  DFFRX1 \R_reg[25][25]  ( .D(n1806), .CK(clk), .RN(reset_n), .Q(\R[25][25] ), 
        .QN(n772) );
  DFFRX1 \R_reg[25][26]  ( .D(n1805), .CK(clk), .RN(reset_n), .Q(\R[25][26] ), 
        .QN(n771) );
  DFFRX1 \R_reg[25][27]  ( .D(n1804), .CK(clk), .RN(reset_n), .Q(\R[25][27] ), 
        .QN(n770) );
  DFFRX1 \R_reg[25][28]  ( .D(n1803), .CK(clk), .RN(reset_n), .Q(\R[25][28] ), 
        .QN(n769) );
  DFFRX1 \R_reg[25][29]  ( .D(n1802), .CK(clk), .RN(reset_n), .Q(\R[25][29] ), 
        .QN(n768) );
  DFFRX1 \R_reg[25][30]  ( .D(n1801), .CK(clk), .RN(reset_n), .Q(\R[25][30] ), 
        .QN(n767) );
  DFFRX1 \R_reg[25][31]  ( .D(n1800), .CK(clk), .RN(reset_n), .Q(\R[25][31] ), 
        .QN(n766) );
  DFFRX1 \R_reg[29][24]  ( .D(n1679), .CK(clk), .RN(reset_n), .Q(\R[29][24] ), 
        .QN(n645) );
  DFFRX1 \R_reg[29][25]  ( .D(n1678), .CK(clk), .RN(reset_n), .Q(\R[29][25] ), 
        .QN(n644) );
  DFFRX1 \R_reg[29][26]  ( .D(n1677), .CK(clk), .RN(reset_n), .Q(\R[29][26] ), 
        .QN(n643) );
  DFFRX1 \R_reg[29][27]  ( .D(n1676), .CK(clk), .RN(reset_n), .Q(\R[29][27] ), 
        .QN(n642) );
  DFFRX1 \R_reg[29][28]  ( .D(n1675), .CK(clk), .RN(reset_n), .Q(\R[29][28] ), 
        .QN(n641) );
  DFFRX1 \R_reg[29][29]  ( .D(n1674), .CK(clk), .RN(reset_n), .Q(\R[29][29] ), 
        .QN(n640) );
  DFFRX1 \R_reg[29][30]  ( .D(n1673), .CK(clk), .RN(reset_n), .Q(\R[29][30] ), 
        .QN(n639) );
  DFFRX1 \R_reg[29][31]  ( .D(n1672), .CK(clk), .RN(reset_n), .Q(\R[29][31] ), 
        .QN(n638) );
  DFFRX1 \R_reg[4][24]  ( .D(n2479), .CK(clk), .RN(reset_n), .Q(\R[4][24] ), 
        .QN(n1445) );
  DFFRX1 \R_reg[4][25]  ( .D(n2478), .CK(clk), .RN(reset_n), .Q(\R[4][25] ), 
        .QN(n1444) );
  DFFRX1 \R_reg[4][26]  ( .D(n2477), .CK(clk), .RN(reset_n), .Q(\R[4][26] ), 
        .QN(n1443) );
  DFFRX1 \R_reg[4][27]  ( .D(n2476), .CK(clk), .RN(reset_n), .Q(\R[4][27] ), 
        .QN(n1442) );
  DFFRX1 \R_reg[4][28]  ( .D(n2475), .CK(clk), .RN(reset_n), .Q(\R[4][28] ), 
        .QN(n1441) );
  DFFRX1 \R_reg[4][29]  ( .D(n2474), .CK(clk), .RN(reset_n), .Q(\R[4][29] ), 
        .QN(n1440) );
  DFFRX1 \R_reg[4][30]  ( .D(n2473), .CK(clk), .RN(reset_n), .Q(\R[4][30] ), 
        .QN(n1439) );
  DFFRX1 \R_reg[4][31]  ( .D(n2472), .CK(clk), .RN(reset_n), .Q(\R[4][31] ), 
        .QN(n1438) );
  DFFRX1 \R_reg[8][24]  ( .D(n2351), .CK(clk), .RN(reset_n), .Q(\R[8][24] ), 
        .QN(n1317) );
  DFFRX1 \R_reg[8][25]  ( .D(n2350), .CK(clk), .RN(reset_n), .Q(\R[8][25] ), 
        .QN(n1316) );
  DFFRX1 \R_reg[8][26]  ( .D(n2349), .CK(clk), .RN(reset_n), .Q(\R[8][26] ), 
        .QN(n1315) );
  DFFRX1 \R_reg[8][27]  ( .D(n2348), .CK(clk), .RN(reset_n), .Q(\R[8][27] ), 
        .QN(n1314) );
  DFFRX1 \R_reg[8][28]  ( .D(n2347), .CK(clk), .RN(reset_n), .Q(\R[8][28] ), 
        .QN(n1313) );
  DFFRX1 \R_reg[8][29]  ( .D(n2346), .CK(clk), .RN(reset_n), .Q(\R[8][29] ), 
        .QN(n1312) );
  DFFRX1 \R_reg[8][30]  ( .D(n2345), .CK(clk), .RN(reset_n), .Q(\R[8][30] ), 
        .QN(n1311) );
  DFFRX1 \R_reg[8][31]  ( .D(n2344), .CK(clk), .RN(reset_n), .Q(\R[8][31] ), 
        .QN(n1310) );
  DFFRX1 \R_reg[12][24]  ( .D(n2223), .CK(clk), .RN(reset_n), .Q(\R[12][24] ), 
        .QN(n1189) );
  DFFRX1 \R_reg[12][25]  ( .D(n2222), .CK(clk), .RN(reset_n), .Q(\R[12][25] ), 
        .QN(n1188) );
  DFFRX1 \R_reg[12][26]  ( .D(n2221), .CK(clk), .RN(reset_n), .Q(\R[12][26] ), 
        .QN(n1187) );
  DFFRX1 \R_reg[12][27]  ( .D(n2220), .CK(clk), .RN(reset_n), .Q(\R[12][27] ), 
        .QN(n1186) );
  DFFRX1 \R_reg[12][28]  ( .D(n2219), .CK(clk), .RN(reset_n), .Q(\R[12][28] ), 
        .QN(n1185) );
  DFFRX1 \R_reg[12][29]  ( .D(n2218), .CK(clk), .RN(reset_n), .Q(\R[12][29] ), 
        .QN(n1184) );
  DFFRX1 \R_reg[12][30]  ( .D(n2217), .CK(clk), .RN(reset_n), .Q(\R[12][30] ), 
        .QN(n1183) );
  DFFRX1 \R_reg[12][31]  ( .D(n2216), .CK(clk), .RN(reset_n), .Q(\R[12][31] ), 
        .QN(n1182) );
  DFFRX1 \R_reg[16][24]  ( .D(n2095), .CK(clk), .RN(reset_n), .Q(\R[16][24] ), 
        .QN(n1061) );
  DFFRX1 \R_reg[16][25]  ( .D(n2094), .CK(clk), .RN(reset_n), .Q(\R[16][25] ), 
        .QN(n1060) );
  DFFRX1 \R_reg[16][26]  ( .D(n2093), .CK(clk), .RN(reset_n), .Q(\R[16][26] ), 
        .QN(n1059) );
  DFFRX1 \R_reg[16][27]  ( .D(n2092), .CK(clk), .RN(reset_n), .Q(\R[16][27] ), 
        .QN(n1058) );
  DFFRX1 \R_reg[16][28]  ( .D(n2091), .CK(clk), .RN(reset_n), .Q(\R[16][28] ), 
        .QN(n1057) );
  DFFRX1 \R_reg[16][29]  ( .D(n2090), .CK(clk), .RN(reset_n), .Q(\R[16][29] ), 
        .QN(n1056) );
  DFFRX1 \R_reg[16][30]  ( .D(n2089), .CK(clk), .RN(reset_n), .Q(\R[16][30] ), 
        .QN(n1055) );
  DFFRX1 \R_reg[16][31]  ( .D(n2088), .CK(clk), .RN(reset_n), .Q(\R[16][31] ), 
        .QN(n1054) );
  DFFRX1 \R_reg[20][24]  ( .D(n1967), .CK(clk), .RN(reset_n), .Q(\R[20][24] ), 
        .QN(n933) );
  DFFRX1 \R_reg[20][25]  ( .D(n1966), .CK(clk), .RN(reset_n), .Q(\R[20][25] ), 
        .QN(n932) );
  DFFRX1 \R_reg[20][26]  ( .D(n1965), .CK(clk), .RN(reset_n), .Q(\R[20][26] ), 
        .QN(n931) );
  DFFRX1 \R_reg[20][27]  ( .D(n1964), .CK(clk), .RN(reset_n), .Q(\R[20][27] ), 
        .QN(n930) );
  DFFRX1 \R_reg[20][28]  ( .D(n1963), .CK(clk), .RN(reset_n), .Q(\R[20][28] ), 
        .QN(n929) );
  DFFRX1 \R_reg[20][29]  ( .D(n1962), .CK(clk), .RN(reset_n), .Q(\R[20][29] ), 
        .QN(n928) );
  DFFRX1 \R_reg[20][30]  ( .D(n1961), .CK(clk), .RN(reset_n), .Q(\R[20][30] ), 
        .QN(n927) );
  DFFRX1 \R_reg[20][31]  ( .D(n1960), .CK(clk), .RN(reset_n), .Q(\R[20][31] ), 
        .QN(n926) );
  DFFRX1 \R_reg[24][24]  ( .D(n1839), .CK(clk), .RN(reset_n), .Q(\R[24][24] ), 
        .QN(n805) );
  DFFRX1 \R_reg[24][25]  ( .D(n1838), .CK(clk), .RN(reset_n), .Q(\R[24][25] ), 
        .QN(n804) );
  DFFRX1 \R_reg[24][26]  ( .D(n1837), .CK(clk), .RN(reset_n), .Q(\R[24][26] ), 
        .QN(n803) );
  DFFRX1 \R_reg[24][27]  ( .D(n1836), .CK(clk), .RN(reset_n), .Q(\R[24][27] ), 
        .QN(n802) );
  DFFRX1 \R_reg[24][28]  ( .D(n1835), .CK(clk), .RN(reset_n), .Q(\R[24][28] ), 
        .QN(n801) );
  DFFRX1 \R_reg[24][29]  ( .D(n1834), .CK(clk), .RN(reset_n), .Q(\R[24][29] ), 
        .QN(n800) );
  DFFRX1 \R_reg[24][30]  ( .D(n1833), .CK(clk), .RN(reset_n), .Q(\R[24][30] ), 
        .QN(n799) );
  DFFRX1 \R_reg[24][31]  ( .D(n1832), .CK(clk), .RN(reset_n), .Q(\R[24][31] ), 
        .QN(n798) );
  DFFRX1 \R_reg[28][24]  ( .D(n1711), .CK(clk), .RN(reset_n), .Q(\R[28][24] ), 
        .QN(n677) );
  DFFRX1 \R_reg[28][25]  ( .D(n1710), .CK(clk), .RN(reset_n), .Q(\R[28][25] ), 
        .QN(n676) );
  DFFRX1 \R_reg[28][26]  ( .D(n1709), .CK(clk), .RN(reset_n), .Q(\R[28][26] ), 
        .QN(n675) );
  DFFRX1 \R_reg[28][27]  ( .D(n1708), .CK(clk), .RN(reset_n), .Q(\R[28][27] ), 
        .QN(n674) );
  DFFRX1 \R_reg[28][28]  ( .D(n1707), .CK(clk), .RN(reset_n), .Q(\R[28][28] ), 
        .QN(n673) );
  DFFRX1 \R_reg[28][29]  ( .D(n1706), .CK(clk), .RN(reset_n), .Q(\R[28][29] ), 
        .QN(n672) );
  DFFRX1 \R_reg[28][30]  ( .D(n1705), .CK(clk), .RN(reset_n), .Q(\R[28][30] ), 
        .QN(n671) );
  DFFRX1 \R_reg[28][31]  ( .D(n1704), .CK(clk), .RN(reset_n), .Q(\R[28][31] ), 
        .QN(n670) );
  DFFRX1 \R_reg[6][24]  ( .D(n2415), .CK(clk), .RN(reset_n), .Q(\R[6][24] ), 
        .QN(n1381) );
  DFFRX1 \R_reg[6][25]  ( .D(n2414), .CK(clk), .RN(reset_n), .Q(\R[6][25] ), 
        .QN(n1380) );
  DFFRX1 \R_reg[6][26]  ( .D(n2413), .CK(clk), .RN(reset_n), .Q(\R[6][26] ), 
        .QN(n1379) );
  DFFRX1 \R_reg[6][27]  ( .D(n2412), .CK(clk), .RN(reset_n), .Q(\R[6][27] ), 
        .QN(n1378) );
  DFFRX1 \R_reg[6][28]  ( .D(n2411), .CK(clk), .RN(reset_n), .Q(\R[6][28] ), 
        .QN(n1377) );
  DFFRX1 \R_reg[6][29]  ( .D(n2410), .CK(clk), .RN(reset_n), .Q(\R[6][29] ), 
        .QN(n1376) );
  DFFRX1 \R_reg[6][30]  ( .D(n2409), .CK(clk), .RN(reset_n), .Q(\R[6][30] ), 
        .QN(n1375) );
  DFFRX1 \R_reg[6][31]  ( .D(n2408), .CK(clk), .RN(reset_n), .Q(\R[6][31] ), 
        .QN(n1374) );
  DFFRX1 \R_reg[10][24]  ( .D(n2287), .CK(clk), .RN(reset_n), .Q(\R[10][24] ), 
        .QN(n1253) );
  DFFRX1 \R_reg[10][25]  ( .D(n2286), .CK(clk), .RN(reset_n), .Q(\R[10][25] ), 
        .QN(n1252) );
  DFFRX1 \R_reg[10][26]  ( .D(n2285), .CK(clk), .RN(reset_n), .Q(\R[10][26] ), 
        .QN(n1251) );
  DFFRX1 \R_reg[10][27]  ( .D(n2284), .CK(clk), .RN(reset_n), .Q(\R[10][27] ), 
        .QN(n1250) );
  DFFRX1 \R_reg[10][28]  ( .D(n2283), .CK(clk), .RN(reset_n), .Q(\R[10][28] ), 
        .QN(n1249) );
  DFFRX1 \R_reg[10][29]  ( .D(n2282), .CK(clk), .RN(reset_n), .Q(\R[10][29] ), 
        .QN(n1248) );
  DFFRX1 \R_reg[10][30]  ( .D(n2281), .CK(clk), .RN(reset_n), .Q(\R[10][30] ), 
        .QN(n1247) );
  DFFRX1 \R_reg[14][24]  ( .D(n2159), .CK(clk), .RN(reset_n), .Q(\R[14][24] ), 
        .QN(n1125) );
  DFFRX1 \R_reg[14][25]  ( .D(n2158), .CK(clk), .RN(reset_n), .Q(\R[14][25] ), 
        .QN(n1124) );
  DFFRX1 \R_reg[14][26]  ( .D(n2157), .CK(clk), .RN(reset_n), .Q(\R[14][26] ), 
        .QN(n1123) );
  DFFRX1 \R_reg[14][27]  ( .D(n2156), .CK(clk), .RN(reset_n), .Q(\R[14][27] ), 
        .QN(n1122) );
  DFFRX1 \R_reg[14][28]  ( .D(n2155), .CK(clk), .RN(reset_n), .Q(\R[14][28] ), 
        .QN(n1121) );
  DFFRX1 \R_reg[14][29]  ( .D(n2154), .CK(clk), .RN(reset_n), .Q(\R[14][29] ), 
        .QN(n1120) );
  DFFRX1 \R_reg[14][30]  ( .D(n2153), .CK(clk), .RN(reset_n), .Q(\R[14][30] ), 
        .QN(n1119) );
  DFFRX1 \R_reg[14][31]  ( .D(n2152), .CK(clk), .RN(reset_n), .Q(\R[14][31] ), 
        .QN(n1118) );
  DFFRX1 \R_reg[18][24]  ( .D(n2031), .CK(clk), .RN(reset_n), .Q(\R[18][24] ), 
        .QN(n997) );
  DFFRX1 \R_reg[18][25]  ( .D(n2030), .CK(clk), .RN(reset_n), .Q(\R[18][25] ), 
        .QN(n996) );
  DFFRX1 \R_reg[18][26]  ( .D(n2029), .CK(clk), .RN(reset_n), .Q(\R[18][26] ), 
        .QN(n995) );
  DFFRX1 \R_reg[18][27]  ( .D(n2028), .CK(clk), .RN(reset_n), .Q(\R[18][27] ), 
        .QN(n994) );
  DFFRX1 \R_reg[18][28]  ( .D(n2027), .CK(clk), .RN(reset_n), .Q(\R[18][28] ), 
        .QN(n993) );
  DFFRX1 \R_reg[18][29]  ( .D(n2026), .CK(clk), .RN(reset_n), .Q(\R[18][29] ), 
        .QN(n992) );
  DFFRX1 \R_reg[18][30]  ( .D(n2025), .CK(clk), .RN(reset_n), .Q(\R[18][30] ), 
        .QN(n991) );
  DFFRX1 \R_reg[18][31]  ( .D(n2024), .CK(clk), .RN(reset_n), .Q(\R[18][31] ), 
        .QN(n990) );
  DFFRX1 \R_reg[22][24]  ( .D(n1903), .CK(clk), .RN(reset_n), .Q(\R[22][24] ), 
        .QN(n869) );
  DFFRX1 \R_reg[22][25]  ( .D(n1902), .CK(clk), .RN(reset_n), .Q(\R[22][25] ), 
        .QN(n868) );
  DFFRX1 \R_reg[22][26]  ( .D(n1901), .CK(clk), .RN(reset_n), .Q(\R[22][26] ), 
        .QN(n867) );
  DFFRX1 \R_reg[22][27]  ( .D(n1900), .CK(clk), .RN(reset_n), .Q(\R[22][27] ), 
        .QN(n866) );
  DFFRX1 \R_reg[22][28]  ( .D(n1899), .CK(clk), .RN(reset_n), .Q(\R[22][28] ), 
        .QN(n865) );
  DFFRX1 \R_reg[22][29]  ( .D(n1898), .CK(clk), .RN(reset_n), .Q(\R[22][29] ), 
        .QN(n864) );
  DFFRX1 \R_reg[22][30]  ( .D(n1897), .CK(clk), .RN(reset_n), .Q(\R[22][30] ), 
        .QN(n863) );
  DFFRX1 \R_reg[22][31]  ( .D(n1896), .CK(clk), .RN(reset_n), .Q(\R[22][31] ), 
        .QN(n862) );
  DFFRX1 \R_reg[26][24]  ( .D(n1775), .CK(clk), .RN(reset_n), .Q(\R[26][24] ), 
        .QN(n741) );
  DFFRX1 \R_reg[26][25]  ( .D(n1774), .CK(clk), .RN(reset_n), .Q(\R[26][25] ), 
        .QN(n740) );
  DFFRX1 \R_reg[26][26]  ( .D(n1773), .CK(clk), .RN(reset_n), .Q(\R[26][26] ), 
        .QN(n739) );
  DFFRX1 \R_reg[26][27]  ( .D(n1772), .CK(clk), .RN(reset_n), .Q(\R[26][27] ), 
        .QN(n738) );
  DFFRX1 \R_reg[26][28]  ( .D(n1771), .CK(clk), .RN(reset_n), .Q(\R[26][28] ), 
        .QN(n737) );
  DFFRX1 \R_reg[26][29]  ( .D(n1770), .CK(clk), .RN(reset_n), .Q(\R[26][29] ), 
        .QN(n736) );
  DFFRX1 \R_reg[26][30]  ( .D(n1769), .CK(clk), .RN(reset_n), .Q(\R[26][30] ), 
        .QN(n735) );
  DFFRX1 \R_reg[26][31]  ( .D(n1768), .CK(clk), .RN(reset_n), .Q(\R[26][31] ), 
        .QN(n734) );
  DFFRX1 \R_reg[30][24]  ( .D(n1647), .CK(clk), .RN(reset_n), .Q(\R[30][24] ), 
        .QN(n613) );
  DFFRX1 \R_reg[30][25]  ( .D(n1646), .CK(clk), .RN(reset_n), .Q(\R[30][25] ), 
        .QN(n612) );
  DFFRX1 \R_reg[30][26]  ( .D(n1645), .CK(clk), .RN(reset_n), .Q(\R[30][26] ), 
        .QN(n611) );
  DFFRX1 \R_reg[30][27]  ( .D(n1644), .CK(clk), .RN(reset_n), .Q(\R[30][27] ), 
        .QN(n610) );
  DFFRX1 \R_reg[30][28]  ( .D(n1643), .CK(clk), .RN(reset_n), .Q(\R[30][28] ), 
        .QN(n609) );
  DFFRX1 \R_reg[30][29]  ( .D(n1642), .CK(clk), .RN(reset_n), .Q(\R[30][29] ), 
        .QN(n608) );
  DFFRX1 \R_reg[30][30]  ( .D(n1641), .CK(clk), .RN(reset_n), .Q(\R[30][30] ), 
        .QN(n607) );
  DFFRX1 \R_reg[30][31]  ( .D(n1640), .CK(clk), .RN(reset_n), .Q(\R[30][31] ), 
        .QN(n606) );
  DFFRX1 \counter_reg[10]  ( .D(N136), .CK(clk), .RN(reset_n), .Q(counter[10]), 
        .QN(n53) );
  DFFRX1 \counter_reg[12]  ( .D(N138), .CK(clk), .RN(reset_n), .Q(counter[12]), 
        .QN(n51) );
  DFFRX1 \counter_reg[11]  ( .D(N137), .CK(clk), .RN(reset_n), .Q(counter[11]), 
        .QN(n52) );
  DFFRX1 \counter_reg[14]  ( .D(N140), .CK(clk), .RN(reset_n), .Q(counter[14]), 
        .QN(n49) );
  DFFRX1 \counter_reg[13]  ( .D(N139), .CK(clk), .RN(reset_n), .Q(counter[13]), 
        .QN(n50) );
  DFFRX1 \counter_reg[15]  ( .D(N141), .CK(clk), .RN(reset_n), .Q(counter[15]), 
        .QN(n48) );
  DFFRX1 \counter_reg[9]  ( .D(N135), .CK(clk), .RN(reset_n), .Q(counter[9]), 
        .QN(n54) );
  DFFRX1 \PC_reg[17]  ( .D(n2612), .CK(clk), .RN(reset_n), .Q(PC[17]), .QN(
        n1578) );
  DFFRX1 \PC_reg[18]  ( .D(n2611), .CK(clk), .RN(reset_n), .Q(PC[18]), .QN(
        n1577) );
  DFFRX1 \PC_reg[19]  ( .D(n2610), .CK(clk), .RN(reset_n), .Q(PC[19]), .QN(
        n1576) );
  DFFRX1 \PC_reg[20]  ( .D(n2609), .CK(clk), .RN(reset_n), .Q(PC[20]), .QN(
        n1575) );
  DFFRX1 \PC_reg[21]  ( .D(n2608), .CK(clk), .RN(reset_n), .Q(PC[21]), .QN(
        n1574) );
  DFFRX1 \R_reg[1][24]  ( .D(n2575), .CK(clk), .RN(reset_n), .Q(\R[1][24] ), 
        .QN(n1541) );
  DFFRX1 \R_reg[1][25]  ( .D(n2574), .CK(clk), .RN(reset_n), .Q(\R[1][25] ), 
        .QN(n1540) );
  DFFRX1 \R_reg[1][26]  ( .D(n2573), .CK(clk), .RN(reset_n), .Q(\R[1][26] ), 
        .QN(n1539) );
  DFFRX1 \R_reg[1][27]  ( .D(n2572), .CK(clk), .RN(reset_n), .Q(\R[1][27] ), 
        .QN(n1538) );
  DFFRX1 \R_reg[1][28]  ( .D(n2571), .CK(clk), .RN(reset_n), .Q(\R[1][28] ), 
        .QN(n1537) );
  DFFRX1 \R_reg[1][29]  ( .D(n2570), .CK(clk), .RN(reset_n), .Q(\R[1][29] ), 
        .QN(n1536) );
  DFFRX1 \R_reg[1][30]  ( .D(n2569), .CK(clk), .RN(reset_n), .Q(\R[1][30] ), 
        .QN(n1535) );
  DFFRX1 \R_reg[1][31]  ( .D(n2568), .CK(clk), .RN(reset_n), .Q(\R[1][31] ), 
        .QN(n1534) );
  DFFRX1 \R_reg[3][24]  ( .D(n2511), .CK(clk), .RN(reset_n), .Q(\R[3][24] ), 
        .QN(n1477) );
  DFFRX1 \R_reg[3][25]  ( .D(n2510), .CK(clk), .RN(reset_n), .Q(\R[3][25] ), 
        .QN(n1476) );
  DFFRX1 \R_reg[3][26]  ( .D(n2509), .CK(clk), .RN(reset_n), .Q(\R[3][26] ), 
        .QN(n1475) );
  DFFRX1 \R_reg[3][27]  ( .D(n2508), .CK(clk), .RN(reset_n), .Q(\R[3][27] ), 
        .QN(n1474) );
  DFFRX1 \R_reg[3][28]  ( .D(n2507), .CK(clk), .RN(reset_n), .Q(\R[3][28] ), 
        .QN(n1473) );
  DFFRX1 \R_reg[3][29]  ( .D(n2506), .CK(clk), .RN(reset_n), .Q(\R[3][29] ), 
        .QN(n1472) );
  DFFRX1 \R_reg[3][30]  ( .D(n2505), .CK(clk), .RN(reset_n), .Q(\R[3][30] ), 
        .QN(n1471) );
  DFFRX1 \R_reg[3][31]  ( .D(n2504), .CK(clk), .RN(reset_n), .Q(\R[3][31] ), 
        .QN(n1470) );
  DFFRX1 \R_reg[2][24]  ( .D(n2543), .CK(clk), .RN(reset_n), .QN(n1509) );
  DFFRX1 \R_reg[2][25]  ( .D(n2542), .CK(clk), .RN(reset_n), .QN(n1508) );
  DFFRX1 \R_reg[2][26]  ( .D(n2541), .CK(clk), .RN(reset_n), .QN(n1507) );
  DFFRX1 \R_reg[2][27]  ( .D(n2540), .CK(clk), .RN(reset_n), .QN(n1506) );
  DFFRX1 \R_reg[2][28]  ( .D(n2539), .CK(clk), .RN(reset_n), .QN(n1505) );
  DFFRX1 \R_reg[2][29]  ( .D(n2538), .CK(clk), .RN(reset_n), .QN(n1504) );
  DFFRX1 \R_reg[2][30]  ( .D(n2537), .CK(clk), .RN(reset_n), .QN(n1503) );
  DFFRX1 \R_reg[2][31]  ( .D(n2536), .CK(clk), .RN(reset_n), .QN(n1502) );
  DFFRX1 \R_reg[7][18]  ( .D(n2389), .CK(clk), .RN(reset_n), .Q(\R[7][18] ), 
        .QN(n1355) );
  DFFRX1 \R_reg[7][19]  ( .D(n2388), .CK(clk), .RN(reset_n), .Q(\R[7][19] ), 
        .QN(n1354) );
  DFFRX1 \R_reg[7][20]  ( .D(n2387), .CK(clk), .RN(reset_n), .Q(\R[7][20] ), 
        .QN(n1353) );
  DFFRX1 \R_reg[7][21]  ( .D(n2386), .CK(clk), .RN(reset_n), .Q(\R[7][21] ), 
        .QN(n1352) );
  DFFRX1 \R_reg[7][22]  ( .D(n2385), .CK(clk), .RN(reset_n), .Q(\R[7][22] ), 
        .QN(n1351) );
  DFFRX1 \R_reg[7][23]  ( .D(n2384), .CK(clk), .RN(reset_n), .Q(\R[7][23] ), 
        .QN(n1350) );
  DFFRX1 \R_reg[11][18]  ( .D(n2261), .CK(clk), .RN(reset_n), .Q(\R[11][18] ), 
        .QN(n1227) );
  DFFRX1 \R_reg[11][19]  ( .D(n2260), .CK(clk), .RN(reset_n), .Q(\R[11][19] ), 
        .QN(n1226) );
  DFFRX1 \R_reg[11][20]  ( .D(n2259), .CK(clk), .RN(reset_n), .Q(\R[11][20] ), 
        .QN(n1225) );
  DFFRX1 \R_reg[11][21]  ( .D(n2258), .CK(clk), .RN(reset_n), .Q(\R[11][21] ), 
        .QN(n1224) );
  DFFRX1 \R_reg[11][22]  ( .D(n2257), .CK(clk), .RN(reset_n), .Q(\R[11][22] ), 
        .QN(n1223) );
  DFFRX1 \R_reg[11][23]  ( .D(n2256), .CK(clk), .RN(reset_n), .Q(\R[11][23] ), 
        .QN(n1222) );
  DFFRX1 \R_reg[15][18]  ( .D(n2133), .CK(clk), .RN(reset_n), .Q(\R[15][18] ), 
        .QN(n1099) );
  DFFRX1 \R_reg[15][19]  ( .D(n2132), .CK(clk), .RN(reset_n), .Q(\R[15][19] ), 
        .QN(n1098) );
  DFFRX1 \R_reg[15][20]  ( .D(n2131), .CK(clk), .RN(reset_n), .Q(\R[15][20] ), 
        .QN(n1097) );
  DFFRX1 \R_reg[15][21]  ( .D(n2130), .CK(clk), .RN(reset_n), .Q(\R[15][21] ), 
        .QN(n1096) );
  DFFRX1 \R_reg[15][22]  ( .D(n2129), .CK(clk), .RN(reset_n), .Q(\R[15][22] ), 
        .QN(n1095) );
  DFFRX1 \R_reg[15][23]  ( .D(n2128), .CK(clk), .RN(reset_n), .Q(\R[15][23] ), 
        .QN(n1094) );
  DFFRX1 \R_reg[19][18]  ( .D(n2005), .CK(clk), .RN(reset_n), .Q(\R[19][18] ), 
        .QN(n971) );
  DFFRX1 \R_reg[19][19]  ( .D(n2004), .CK(clk), .RN(reset_n), .Q(\R[19][19] ), 
        .QN(n970) );
  DFFRX1 \R_reg[19][20]  ( .D(n2003), .CK(clk), .RN(reset_n), .Q(\R[19][20] ), 
        .QN(n969) );
  DFFRX1 \R_reg[19][21]  ( .D(n2002), .CK(clk), .RN(reset_n), .Q(\R[19][21] ), 
        .QN(n968) );
  DFFRX1 \R_reg[19][22]  ( .D(n2001), .CK(clk), .RN(reset_n), .Q(\R[19][22] ), 
        .QN(n967) );
  DFFRX1 \R_reg[19][23]  ( .D(n2000), .CK(clk), .RN(reset_n), .Q(\R[19][23] ), 
        .QN(n966) );
  DFFRX1 \R_reg[23][18]  ( .D(n1877), .CK(clk), .RN(reset_n), .Q(\R[23][18] ), 
        .QN(n843) );
  DFFRX1 \R_reg[23][19]  ( .D(n1876), .CK(clk), .RN(reset_n), .Q(\R[23][19] ), 
        .QN(n842) );
  DFFRX1 \R_reg[23][20]  ( .D(n1875), .CK(clk), .RN(reset_n), .Q(\R[23][20] ), 
        .QN(n841) );
  DFFRX1 \R_reg[23][21]  ( .D(n1874), .CK(clk), .RN(reset_n), .Q(\R[23][21] ), 
        .QN(n840) );
  DFFRX1 \R_reg[23][22]  ( .D(n1873), .CK(clk), .RN(reset_n), .Q(\R[23][22] ), 
        .QN(n839) );
  DFFRX1 \R_reg[23][23]  ( .D(n1872), .CK(clk), .RN(reset_n), .Q(\R[23][23] ), 
        .QN(n838) );
  DFFRX1 \R_reg[27][18]  ( .D(n1749), .CK(clk), .RN(reset_n), .Q(\R[27][18] ), 
        .QN(n715) );
  DFFRX1 \R_reg[27][19]  ( .D(n1748), .CK(clk), .RN(reset_n), .Q(\R[27][19] ), 
        .QN(n714) );
  DFFRX1 \R_reg[27][20]  ( .D(n1747), .CK(clk), .RN(reset_n), .Q(\R[27][20] ), 
        .QN(n713) );
  DFFRX1 \R_reg[27][21]  ( .D(n1746), .CK(clk), .RN(reset_n), .Q(\R[27][21] ), 
        .QN(n712) );
  DFFRX1 \R_reg[27][22]  ( .D(n1745), .CK(clk), .RN(reset_n), .Q(\R[27][22] ), 
        .QN(n711) );
  DFFRX1 \R_reg[27][23]  ( .D(n1744), .CK(clk), .RN(reset_n), .Q(\R[27][23] ), 
        .QN(n710) );
  DFFRX1 \R_reg[31][18]  ( .D(n1621), .CK(clk), .RN(reset_n), .Q(\R[31][18] ), 
        .QN(n587) );
  DFFRX1 \R_reg[31][19]  ( .D(n1620), .CK(clk), .RN(reset_n), .Q(\R[31][19] ), 
        .QN(n586) );
  DFFRX1 \R_reg[31][20]  ( .D(n1619), .CK(clk), .RN(reset_n), .Q(\R[31][20] ), 
        .QN(n585) );
  DFFRX1 \R_reg[31][21]  ( .D(n1618), .CK(clk), .RN(reset_n), .Q(\R[31][21] ), 
        .QN(n584) );
  DFFRX1 \R_reg[31][22]  ( .D(n1617), .CK(clk), .RN(reset_n), .Q(\R[31][22] ), 
        .QN(n583) );
  DFFRX1 \R_reg[31][23]  ( .D(n1616), .CK(clk), .RN(reset_n), .Q(\R[31][23] ), 
        .QN(n582) );
  DFFRX1 \R_reg[5][18]  ( .D(n2453), .CK(clk), .RN(reset_n), .Q(\R[5][18] ), 
        .QN(n1419) );
  DFFRX1 \R_reg[5][19]  ( .D(n2452), .CK(clk), .RN(reset_n), .Q(\R[5][19] ), 
        .QN(n1418) );
  DFFRX1 \R_reg[5][20]  ( .D(n2451), .CK(clk), .RN(reset_n), .Q(\R[5][20] ), 
        .QN(n1417) );
  DFFRX1 \R_reg[5][21]  ( .D(n2450), .CK(clk), .RN(reset_n), .Q(\R[5][21] ), 
        .QN(n1416) );
  DFFRX1 \R_reg[5][22]  ( .D(n2449), .CK(clk), .RN(reset_n), .Q(\R[5][22] ), 
        .QN(n1415) );
  DFFRX1 \R_reg[5][23]  ( .D(n2448), .CK(clk), .RN(reset_n), .Q(\R[5][23] ), 
        .QN(n1414) );
  DFFRX1 \R_reg[9][19]  ( .D(n2324), .CK(clk), .RN(reset_n), .Q(\R[9][19] ), 
        .QN(n1290) );
  DFFRX1 \R_reg[9][20]  ( .D(n2323), .CK(clk), .RN(reset_n), .Q(\R[9][20] ), 
        .QN(n1289) );
  DFFRX1 \R_reg[9][21]  ( .D(n2322), .CK(clk), .RN(reset_n), .Q(\R[9][21] ), 
        .QN(n1288) );
  DFFRX1 \R_reg[9][22]  ( .D(n2321), .CK(clk), .RN(reset_n), .Q(\R[9][22] ), 
        .QN(n1287) );
  DFFRX1 \R_reg[9][23]  ( .D(n2320), .CK(clk), .RN(reset_n), .Q(\R[9][23] ), 
        .QN(n1286) );
  DFFRX1 \R_reg[13][18]  ( .D(n2197), .CK(clk), .RN(reset_n), .Q(\R[13][18] ), 
        .QN(n1163) );
  DFFRX1 \R_reg[13][19]  ( .D(n2196), .CK(clk), .RN(reset_n), .Q(\R[13][19] ), 
        .QN(n1162) );
  DFFRX1 \R_reg[13][20]  ( .D(n2195), .CK(clk), .RN(reset_n), .Q(\R[13][20] ), 
        .QN(n1161) );
  DFFRX1 \R_reg[13][21]  ( .D(n2194), .CK(clk), .RN(reset_n), .Q(\R[13][21] ), 
        .QN(n1160) );
  DFFRX1 \R_reg[13][22]  ( .D(n2193), .CK(clk), .RN(reset_n), .Q(\R[13][22] ), 
        .QN(n1159) );
  DFFRX1 \R_reg[13][23]  ( .D(n2192), .CK(clk), .RN(reset_n), .Q(\R[13][23] ), 
        .QN(n1158) );
  DFFRX1 \R_reg[17][19]  ( .D(n2068), .CK(clk), .RN(reset_n), .Q(\R[17][19] ), 
        .QN(n1034) );
  DFFRX1 \R_reg[17][20]  ( .D(n2067), .CK(clk), .RN(reset_n), .Q(\R[17][20] ), 
        .QN(n1033) );
  DFFRX1 \R_reg[17][21]  ( .D(n2066), .CK(clk), .RN(reset_n), .Q(\R[17][21] ), 
        .QN(n1032) );
  DFFRX1 \R_reg[17][22]  ( .D(n2065), .CK(clk), .RN(reset_n), .Q(\R[17][22] ), 
        .QN(n1031) );
  DFFRX1 \R_reg[17][23]  ( .D(n2064), .CK(clk), .RN(reset_n), .Q(\R[17][23] ), 
        .QN(n1030) );
  DFFRX1 \R_reg[21][18]  ( .D(n1941), .CK(clk), .RN(reset_n), .Q(\R[21][18] ), 
        .QN(n907) );
  DFFRX1 \R_reg[21][19]  ( .D(n1940), .CK(clk), .RN(reset_n), .Q(\R[21][19] ), 
        .QN(n906) );
  DFFRX1 \R_reg[21][20]  ( .D(n1939), .CK(clk), .RN(reset_n), .Q(\R[21][20] ), 
        .QN(n905) );
  DFFRX1 \R_reg[21][21]  ( .D(n1938), .CK(clk), .RN(reset_n), .Q(\R[21][21] ), 
        .QN(n904) );
  DFFRX1 \R_reg[21][22]  ( .D(n1937), .CK(clk), .RN(reset_n), .Q(\R[21][22] ), 
        .QN(n903) );
  DFFRX1 \R_reg[21][23]  ( .D(n1936), .CK(clk), .RN(reset_n), .Q(\R[21][23] ), 
        .QN(n902) );
  DFFRX1 \R_reg[25][19]  ( .D(n1812), .CK(clk), .RN(reset_n), .Q(\R[25][19] ), 
        .QN(n778) );
  DFFRX1 \R_reg[25][20]  ( .D(n1811), .CK(clk), .RN(reset_n), .Q(\R[25][20] ), 
        .QN(n777) );
  DFFRX1 \R_reg[25][21]  ( .D(n1810), .CK(clk), .RN(reset_n), .Q(\R[25][21] ), 
        .QN(n776) );
  DFFRX1 \R_reg[25][22]  ( .D(n1809), .CK(clk), .RN(reset_n), .Q(\R[25][22] ), 
        .QN(n775) );
  DFFRX1 \R_reg[25][23]  ( .D(n1808), .CK(clk), .RN(reset_n), .Q(\R[25][23] ), 
        .QN(n774) );
  DFFRX1 \R_reg[29][18]  ( .D(n1685), .CK(clk), .RN(reset_n), .Q(\R[29][18] ), 
        .QN(n651) );
  DFFRX1 \R_reg[29][19]  ( .D(n1684), .CK(clk), .RN(reset_n), .Q(\R[29][19] ), 
        .QN(n650) );
  DFFRX1 \R_reg[29][20]  ( .D(n1683), .CK(clk), .RN(reset_n), .Q(\R[29][20] ), 
        .QN(n649) );
  DFFRX1 \R_reg[29][21]  ( .D(n1682), .CK(clk), .RN(reset_n), .Q(\R[29][21] ), 
        .QN(n648) );
  DFFRX1 \R_reg[29][22]  ( .D(n1681), .CK(clk), .RN(reset_n), .Q(\R[29][22] ), 
        .QN(n647) );
  DFFRX1 \R_reg[29][23]  ( .D(n1680), .CK(clk), .RN(reset_n), .Q(\R[29][23] ), 
        .QN(n646) );
  DFFRX1 \R_reg[4][18]  ( .D(n2485), .CK(clk), .RN(reset_n), .Q(\R[4][18] ), 
        .QN(n1451) );
  DFFRX1 \R_reg[4][19]  ( .D(n2484), .CK(clk), .RN(reset_n), .Q(\R[4][19] ), 
        .QN(n1450) );
  DFFRX1 \R_reg[4][20]  ( .D(n2483), .CK(clk), .RN(reset_n), .Q(\R[4][20] ), 
        .QN(n1449) );
  DFFRX1 \R_reg[4][21]  ( .D(n2482), .CK(clk), .RN(reset_n), .Q(\R[4][21] ), 
        .QN(n1448) );
  DFFRX1 \R_reg[4][22]  ( .D(n2481), .CK(clk), .RN(reset_n), .Q(\R[4][22] ), 
        .QN(n1447) );
  DFFRX1 \R_reg[4][23]  ( .D(n2480), .CK(clk), .RN(reset_n), .Q(\R[4][23] ), 
        .QN(n1446) );
  DFFRX1 \R_reg[8][19]  ( .D(n2356), .CK(clk), .RN(reset_n), .Q(\R[8][19] ), 
        .QN(n1322) );
  DFFRX1 \R_reg[8][20]  ( .D(n2355), .CK(clk), .RN(reset_n), .Q(\R[8][20] ), 
        .QN(n1321) );
  DFFRX1 \R_reg[8][21]  ( .D(n2354), .CK(clk), .RN(reset_n), .Q(\R[8][21] ), 
        .QN(n1320) );
  DFFRX1 \R_reg[8][22]  ( .D(n2353), .CK(clk), .RN(reset_n), .Q(\R[8][22] ), 
        .QN(n1319) );
  DFFRX1 \R_reg[8][23]  ( .D(n2352), .CK(clk), .RN(reset_n), .Q(\R[8][23] ), 
        .QN(n1318) );
  DFFRX1 \R_reg[12][18]  ( .D(n2229), .CK(clk), .RN(reset_n), .Q(\R[12][18] ), 
        .QN(n1195) );
  DFFRX1 \R_reg[12][19]  ( .D(n2228), .CK(clk), .RN(reset_n), .Q(\R[12][19] ), 
        .QN(n1194) );
  DFFRX1 \R_reg[12][20]  ( .D(n2227), .CK(clk), .RN(reset_n), .Q(\R[12][20] ), 
        .QN(n1193) );
  DFFRX1 \R_reg[12][21]  ( .D(n2226), .CK(clk), .RN(reset_n), .Q(\R[12][21] ), 
        .QN(n1192) );
  DFFRX1 \R_reg[12][22]  ( .D(n2225), .CK(clk), .RN(reset_n), .Q(\R[12][22] ), 
        .QN(n1191) );
  DFFRX1 \R_reg[12][23]  ( .D(n2224), .CK(clk), .RN(reset_n), .Q(\R[12][23] ), 
        .QN(n1190) );
  DFFRX1 \R_reg[16][19]  ( .D(n2100), .CK(clk), .RN(reset_n), .Q(\R[16][19] ), 
        .QN(n1066) );
  DFFRX1 \R_reg[16][20]  ( .D(n2099), .CK(clk), .RN(reset_n), .Q(\R[16][20] ), 
        .QN(n1065) );
  DFFRX1 \R_reg[16][21]  ( .D(n2098), .CK(clk), .RN(reset_n), .Q(\R[16][21] ), 
        .QN(n1064) );
  DFFRX1 \R_reg[16][22]  ( .D(n2097), .CK(clk), .RN(reset_n), .Q(\R[16][22] ), 
        .QN(n1063) );
  DFFRX1 \R_reg[16][23]  ( .D(n2096), .CK(clk), .RN(reset_n), .Q(\R[16][23] ), 
        .QN(n1062) );
  DFFRX1 \R_reg[20][18]  ( .D(n1973), .CK(clk), .RN(reset_n), .Q(\R[20][18] ), 
        .QN(n939) );
  DFFRX1 \R_reg[20][19]  ( .D(n1972), .CK(clk), .RN(reset_n), .Q(\R[20][19] ), 
        .QN(n938) );
  DFFRX1 \R_reg[20][20]  ( .D(n1971), .CK(clk), .RN(reset_n), .Q(\R[20][20] ), 
        .QN(n937) );
  DFFRX1 \R_reg[20][21]  ( .D(n1970), .CK(clk), .RN(reset_n), .Q(\R[20][21] ), 
        .QN(n936) );
  DFFRX1 \R_reg[20][22]  ( .D(n1969), .CK(clk), .RN(reset_n), .Q(\R[20][22] ), 
        .QN(n935) );
  DFFRX1 \R_reg[20][23]  ( .D(n1968), .CK(clk), .RN(reset_n), .Q(\R[20][23] ), 
        .QN(n934) );
  DFFRX1 \R_reg[24][19]  ( .D(n1844), .CK(clk), .RN(reset_n), .Q(\R[24][19] ), 
        .QN(n810) );
  DFFRX1 \R_reg[24][20]  ( .D(n1843), .CK(clk), .RN(reset_n), .Q(\R[24][20] ), 
        .QN(n809) );
  DFFRX1 \R_reg[24][21]  ( .D(n1842), .CK(clk), .RN(reset_n), .Q(\R[24][21] ), 
        .QN(n808) );
  DFFRX1 \R_reg[24][22]  ( .D(n1841), .CK(clk), .RN(reset_n), .Q(\R[24][22] ), 
        .QN(n807) );
  DFFRX1 \R_reg[24][23]  ( .D(n1840), .CK(clk), .RN(reset_n), .Q(\R[24][23] ), 
        .QN(n806) );
  DFFRX1 \R_reg[28][18]  ( .D(n1717), .CK(clk), .RN(reset_n), .Q(\R[28][18] ), 
        .QN(n683) );
  DFFRX1 \R_reg[28][19]  ( .D(n1716), .CK(clk), .RN(reset_n), .Q(\R[28][19] ), 
        .QN(n682) );
  DFFRX1 \R_reg[28][20]  ( .D(n1715), .CK(clk), .RN(reset_n), .Q(\R[28][20] ), 
        .QN(n681) );
  DFFRX1 \R_reg[28][21]  ( .D(n1714), .CK(clk), .RN(reset_n), .Q(\R[28][21] ), 
        .QN(n680) );
  DFFRX1 \R_reg[28][22]  ( .D(n1713), .CK(clk), .RN(reset_n), .Q(\R[28][22] ), 
        .QN(n679) );
  DFFRX1 \R_reg[28][23]  ( .D(n1712), .CK(clk), .RN(reset_n), .Q(\R[28][23] ), 
        .QN(n678) );
  DFFRX1 \R_reg[6][18]  ( .D(n2421), .CK(clk), .RN(reset_n), .Q(\R[6][18] ), 
        .QN(n1387) );
  DFFRX1 \R_reg[6][19]  ( .D(n2420), .CK(clk), .RN(reset_n), .Q(\R[6][19] ), 
        .QN(n1386) );
  DFFRX1 \R_reg[6][20]  ( .D(n2419), .CK(clk), .RN(reset_n), .Q(\R[6][20] ), 
        .QN(n1385) );
  DFFRX1 \R_reg[6][21]  ( .D(n2418), .CK(clk), .RN(reset_n), .Q(\R[6][21] ), 
        .QN(n1384) );
  DFFRX1 \R_reg[6][22]  ( .D(n2417), .CK(clk), .RN(reset_n), .Q(\R[6][22] ), 
        .QN(n1383) );
  DFFRX1 \R_reg[6][23]  ( .D(n2416), .CK(clk), .RN(reset_n), .Q(\R[6][23] ), 
        .QN(n1382) );
  DFFRX1 \R_reg[10][18]  ( .D(n2293), .CK(clk), .RN(reset_n), .Q(\R[10][18] ), 
        .QN(n1259) );
  DFFRX1 \R_reg[10][19]  ( .D(n2292), .CK(clk), .RN(reset_n), .Q(\R[10][19] ), 
        .QN(n1258) );
  DFFRX1 \R_reg[10][20]  ( .D(n2291), .CK(clk), .RN(reset_n), .Q(\R[10][20] ), 
        .QN(n1257) );
  DFFRX1 \R_reg[10][21]  ( .D(n2290), .CK(clk), .RN(reset_n), .Q(\R[10][21] ), 
        .QN(n1256) );
  DFFRX1 \R_reg[10][22]  ( .D(n2289), .CK(clk), .RN(reset_n), .Q(\R[10][22] ), 
        .QN(n1255) );
  DFFRX1 \R_reg[10][23]  ( .D(n2288), .CK(clk), .RN(reset_n), .Q(\R[10][23] ), 
        .QN(n1254) );
  DFFRX1 \R_reg[14][18]  ( .D(n2165), .CK(clk), .RN(reset_n), .Q(\R[14][18] ), 
        .QN(n1131) );
  DFFRX1 \R_reg[14][19]  ( .D(n2164), .CK(clk), .RN(reset_n), .Q(\R[14][19] ), 
        .QN(n1130) );
  DFFRX1 \R_reg[14][20]  ( .D(n2163), .CK(clk), .RN(reset_n), .Q(\R[14][20] ), 
        .QN(n1129) );
  DFFRX1 \R_reg[14][21]  ( .D(n2162), .CK(clk), .RN(reset_n), .Q(\R[14][21] ), 
        .QN(n1128) );
  DFFRX1 \R_reg[14][22]  ( .D(n2161), .CK(clk), .RN(reset_n), .Q(\R[14][22] ), 
        .QN(n1127) );
  DFFRX1 \R_reg[14][23]  ( .D(n2160), .CK(clk), .RN(reset_n), .Q(\R[14][23] ), 
        .QN(n1126) );
  DFFRX1 \R_reg[18][18]  ( .D(n2037), .CK(clk), .RN(reset_n), .Q(\R[18][18] ), 
        .QN(n1003) );
  DFFRX1 \R_reg[18][19]  ( .D(n2036), .CK(clk), .RN(reset_n), .Q(\R[18][19] ), 
        .QN(n1002) );
  DFFRX1 \R_reg[18][20]  ( .D(n2035), .CK(clk), .RN(reset_n), .Q(\R[18][20] ), 
        .QN(n1001) );
  DFFRX1 \R_reg[18][21]  ( .D(n2034), .CK(clk), .RN(reset_n), .Q(\R[18][21] ), 
        .QN(n1000) );
  DFFRX1 \R_reg[18][22]  ( .D(n2033), .CK(clk), .RN(reset_n), .Q(\R[18][22] ), 
        .QN(n999) );
  DFFRX1 \R_reg[18][23]  ( .D(n2032), .CK(clk), .RN(reset_n), .Q(\R[18][23] ), 
        .QN(n998) );
  DFFRX1 \R_reg[22][18]  ( .D(n1909), .CK(clk), .RN(reset_n), .Q(\R[22][18] ), 
        .QN(n875) );
  DFFRX1 \R_reg[22][19]  ( .D(n1908), .CK(clk), .RN(reset_n), .Q(\R[22][19] ), 
        .QN(n874) );
  DFFRX1 \R_reg[22][20]  ( .D(n1907), .CK(clk), .RN(reset_n), .Q(\R[22][20] ), 
        .QN(n873) );
  DFFRX1 \R_reg[22][21]  ( .D(n1906), .CK(clk), .RN(reset_n), .Q(\R[22][21] ), 
        .QN(n872) );
  DFFRX1 \R_reg[22][22]  ( .D(n1905), .CK(clk), .RN(reset_n), .Q(\R[22][22] ), 
        .QN(n871) );
  DFFRX1 \R_reg[22][23]  ( .D(n1904), .CK(clk), .RN(reset_n), .Q(\R[22][23] ), 
        .QN(n870) );
  DFFRX1 \R_reg[26][18]  ( .D(n1781), .CK(clk), .RN(reset_n), .Q(\R[26][18] ), 
        .QN(n747) );
  DFFRX1 \R_reg[26][19]  ( .D(n1780), .CK(clk), .RN(reset_n), .Q(\R[26][19] ), 
        .QN(n746) );
  DFFRX1 \R_reg[26][20]  ( .D(n1779), .CK(clk), .RN(reset_n), .Q(\R[26][20] ), 
        .QN(n745) );
  DFFRX1 \R_reg[26][21]  ( .D(n1778), .CK(clk), .RN(reset_n), .Q(\R[26][21] ), 
        .QN(n744) );
  DFFRX1 \R_reg[26][22]  ( .D(n1777), .CK(clk), .RN(reset_n), .Q(\R[26][22] ), 
        .QN(n743) );
  DFFRX1 \R_reg[26][23]  ( .D(n1776), .CK(clk), .RN(reset_n), .Q(\R[26][23] ), 
        .QN(n742) );
  DFFRX1 \R_reg[30][18]  ( .D(n1653), .CK(clk), .RN(reset_n), .Q(\R[30][18] ), 
        .QN(n619) );
  DFFRX1 \R_reg[30][19]  ( .D(n1652), .CK(clk), .RN(reset_n), .Q(\R[30][19] ), 
        .QN(n618) );
  DFFRX1 \R_reg[30][20]  ( .D(n1651), .CK(clk), .RN(reset_n), .Q(\R[30][20] ), 
        .QN(n617) );
  DFFRX1 \R_reg[30][21]  ( .D(n1650), .CK(clk), .RN(reset_n), .Q(\R[30][21] ), 
        .QN(n616) );
  DFFRX1 \R_reg[30][22]  ( .D(n1649), .CK(clk), .RN(reset_n), .Q(\R[30][22] ), 
        .QN(n615) );
  DFFRX1 \R_reg[30][23]  ( .D(n1648), .CK(clk), .RN(reset_n), .Q(\R[30][23] ), 
        .QN(n614) );
  DFFRX1 \counter_reg[6]  ( .D(N132), .CK(clk), .RN(reset_n), .Q(counter[6]), 
        .QN(n57) );
  DFFRX1 \counter_reg[8]  ( .D(N134), .CK(clk), .RN(reset_n), .Q(counter[8]), 
        .QN(n55) );
  DFFRX1 \counter_reg[4]  ( .D(N130), .CK(clk), .RN(reset_n), .Q(counter[4]), 
        .QN(n59) );
  DFFRX1 \counter_reg[2]  ( .D(N128), .CK(clk), .RN(reset_n), .Q(counter[2]), 
        .QN(n61) );
  DFFRX1 \counter_reg[7]  ( .D(N133), .CK(clk), .RN(reset_n), .Q(counter[7]), 
        .QN(n56) );
  DFFRX1 \counter_reg[3]  ( .D(N129), .CK(clk), .RN(reset_n), .Q(counter[3]), 
        .QN(n60) );
  DFFRX1 \counter_reg[5]  ( .D(N131), .CK(clk), .RN(reset_n), .Q(counter[5]), 
        .QN(n58) );
  DFFRX1 \PC_reg[11]  ( .D(n2618), .CK(clk), .RN(reset_n), .Q(PC[11]), .QN(
        n1584) );
  DFFRX1 \PC_reg[12]  ( .D(n2617), .CK(clk), .RN(reset_n), .Q(PC[12]), .QN(
        n1583) );
  DFFRX1 \PC_reg[13]  ( .D(n2616), .CK(clk), .RN(reset_n), .Q(PC[13]), .QN(
        n1582) );
  DFFRX1 \PC_reg[14]  ( .D(n2615), .CK(clk), .RN(reset_n), .Q(PC[14]), .QN(
        n1581) );
  DFFRX1 \PC_reg[15]  ( .D(n2614), .CK(clk), .RN(reset_n), .Q(PC[15]), .QN(
        n1580) );
  DFFRX1 \PC_reg[16]  ( .D(n2613), .CK(clk), .RN(reset_n), .Q(PC[16]), .QN(
        n1579) );
  DFFRX1 \R_reg[1][18]  ( .D(n2581), .CK(clk), .RN(reset_n), .Q(\R[1][18] ), 
        .QN(n1547) );
  DFFRX1 \R_reg[1][19]  ( .D(n2580), .CK(clk), .RN(reset_n), .Q(\R[1][19] ), 
        .QN(n1546) );
  DFFRX1 \R_reg[1][20]  ( .D(n2579), .CK(clk), .RN(reset_n), .Q(\R[1][20] ), 
        .QN(n1545) );
  DFFRX1 \R_reg[1][21]  ( .D(n2578), .CK(clk), .RN(reset_n), .Q(\R[1][21] ), 
        .QN(n1544) );
  DFFRX1 \R_reg[1][22]  ( .D(n2577), .CK(clk), .RN(reset_n), .Q(\R[1][22] ), 
        .QN(n1543) );
  DFFRX1 \R_reg[1][23]  ( .D(n2576), .CK(clk), .RN(reset_n), .Q(\R[1][23] ), 
        .QN(n1542) );
  DFFRX1 \R_reg[3][18]  ( .D(n2517), .CK(clk), .RN(reset_n), .Q(\R[3][18] ), 
        .QN(n1483) );
  DFFRX1 \R_reg[3][19]  ( .D(n2516), .CK(clk), .RN(reset_n), .Q(\R[3][19] ), 
        .QN(n1482) );
  DFFRX1 \R_reg[3][20]  ( .D(n2515), .CK(clk), .RN(reset_n), .Q(\R[3][20] ), 
        .QN(n1481) );
  DFFRX1 \R_reg[3][21]  ( .D(n2514), .CK(clk), .RN(reset_n), .Q(\R[3][21] ), 
        .QN(n1480) );
  DFFRX1 \R_reg[3][22]  ( .D(n2513), .CK(clk), .RN(reset_n), .Q(\R[3][22] ), 
        .QN(n1479) );
  DFFRX1 \R_reg[3][23]  ( .D(n2512), .CK(clk), .RN(reset_n), .Q(\R[3][23] ), 
        .QN(n1478) );
  DFFRX1 \R_reg[2][18]  ( .D(n2549), .CK(clk), .RN(reset_n), .QN(n1515) );
  DFFRX1 \R_reg[2][19]  ( .D(n2548), .CK(clk), .RN(reset_n), .QN(n1514) );
  DFFRX1 \R_reg[2][20]  ( .D(n2547), .CK(clk), .RN(reset_n), .QN(n1513) );
  DFFRX1 \R_reg[2][21]  ( .D(n2546), .CK(clk), .RN(reset_n), .QN(n1512) );
  DFFRX1 \R_reg[2][22]  ( .D(n2545), .CK(clk), .RN(reset_n), .QN(n1511) );
  DFFRX1 \R_reg[2][23]  ( .D(n2544), .CK(clk), .RN(reset_n), .QN(n1510) );
  DFFRX1 \R_reg[7][13]  ( .D(n2394), .CK(clk), .RN(reset_n), .Q(\R[7][13] ), 
        .QN(n1360) );
  DFFRX1 \R_reg[7][14]  ( .D(n2393), .CK(clk), .RN(reset_n), .Q(\R[7][14] ), 
        .QN(n1359) );
  DFFRX1 \R_reg[7][15]  ( .D(n2392), .CK(clk), .RN(reset_n), .Q(\R[7][15] ), 
        .QN(n1358) );
  DFFRX1 \R_reg[7][16]  ( .D(n2391), .CK(clk), .RN(reset_n), .Q(\R[7][16] ), 
        .QN(n1357) );
  DFFRX1 \R_reg[7][17]  ( .D(n2390), .CK(clk), .RN(reset_n), .Q(\R[7][17] ), 
        .QN(n1356) );
  DFFRX1 \R_reg[11][13]  ( .D(n2266), .CK(clk), .RN(reset_n), .Q(\R[11][13] ), 
        .QN(n1232) );
  DFFRX1 \R_reg[11][14]  ( .D(n2265), .CK(clk), .RN(reset_n), .Q(\R[11][14] ), 
        .QN(n1231) );
  DFFRX1 \R_reg[11][15]  ( .D(n2264), .CK(clk), .RN(reset_n), .Q(\R[11][15] ), 
        .QN(n1230) );
  DFFRX1 \R_reg[11][16]  ( .D(n2263), .CK(clk), .RN(reset_n), .Q(\R[11][16] ), 
        .QN(n1229) );
  DFFRX1 \R_reg[11][17]  ( .D(n2262), .CK(clk), .RN(reset_n), .Q(\R[11][17] ), 
        .QN(n1228) );
  DFFRX1 \R_reg[15][13]  ( .D(n2138), .CK(clk), .RN(reset_n), .Q(\R[15][13] ), 
        .QN(n1104) );
  DFFRX1 \R_reg[15][14]  ( .D(n2137), .CK(clk), .RN(reset_n), .Q(\R[15][14] ), 
        .QN(n1103) );
  DFFRX1 \R_reg[15][15]  ( .D(n2136), .CK(clk), .RN(reset_n), .Q(\R[15][15] ), 
        .QN(n1102) );
  DFFRX1 \R_reg[15][16]  ( .D(n2135), .CK(clk), .RN(reset_n), .Q(\R[15][16] ), 
        .QN(n1101) );
  DFFRX1 \R_reg[15][17]  ( .D(n2134), .CK(clk), .RN(reset_n), .Q(\R[15][17] ), 
        .QN(n1100) );
  DFFRX1 \R_reg[19][13]  ( .D(n2010), .CK(clk), .RN(reset_n), .Q(\R[19][13] ), 
        .QN(n976) );
  DFFRX1 \R_reg[19][14]  ( .D(n2009), .CK(clk), .RN(reset_n), .Q(\R[19][14] ), 
        .QN(n975) );
  DFFRX1 \R_reg[19][15]  ( .D(n2008), .CK(clk), .RN(reset_n), .Q(\R[19][15] ), 
        .QN(n974) );
  DFFRX1 \R_reg[19][16]  ( .D(n2007), .CK(clk), .RN(reset_n), .Q(\R[19][16] ), 
        .QN(n973) );
  DFFRX1 \R_reg[19][17]  ( .D(n2006), .CK(clk), .RN(reset_n), .Q(\R[19][17] ), 
        .QN(n972) );
  DFFRX1 \R_reg[23][13]  ( .D(n1882), .CK(clk), .RN(reset_n), .Q(\R[23][13] ), 
        .QN(n848) );
  DFFRX1 \R_reg[23][14]  ( .D(n1881), .CK(clk), .RN(reset_n), .Q(\R[23][14] ), 
        .QN(n847) );
  DFFRX1 \R_reg[23][15]  ( .D(n1880), .CK(clk), .RN(reset_n), .Q(\R[23][15] ), 
        .QN(n846) );
  DFFRX1 \R_reg[23][16]  ( .D(n1879), .CK(clk), .RN(reset_n), .Q(\R[23][16] ), 
        .QN(n845) );
  DFFRX1 \R_reg[23][17]  ( .D(n1878), .CK(clk), .RN(reset_n), .Q(\R[23][17] ), 
        .QN(n844) );
  DFFRX1 \R_reg[27][13]  ( .D(n1754), .CK(clk), .RN(reset_n), .Q(\R[27][13] ), 
        .QN(n720) );
  DFFRX1 \R_reg[27][14]  ( .D(n1753), .CK(clk), .RN(reset_n), .Q(\R[27][14] ), 
        .QN(n719) );
  DFFRX1 \R_reg[27][15]  ( .D(n1752), .CK(clk), .RN(reset_n), .Q(\R[27][15] ), 
        .QN(n718) );
  DFFRX1 \R_reg[27][16]  ( .D(n1751), .CK(clk), .RN(reset_n), .Q(\R[27][16] ), 
        .QN(n717) );
  DFFRX1 \R_reg[27][17]  ( .D(n1750), .CK(clk), .RN(reset_n), .Q(\R[27][17] ), 
        .QN(n716) );
  DFFRX1 \R_reg[31][13]  ( .D(n1626), .CK(clk), .RN(reset_n), .Q(\R[31][13] ), 
        .QN(n592) );
  DFFRX1 \R_reg[31][14]  ( .D(n1625), .CK(clk), .RN(reset_n), .Q(\R[31][14] ), 
        .QN(n591) );
  DFFRX1 \R_reg[31][15]  ( .D(n1624), .CK(clk), .RN(reset_n), .Q(\R[31][15] ), 
        .QN(n590) );
  DFFRX1 \R_reg[31][16]  ( .D(n1623), .CK(clk), .RN(reset_n), .Q(\R[31][16] ), 
        .QN(n589) );
  DFFRX1 \R_reg[31][17]  ( .D(n1622), .CK(clk), .RN(reset_n), .Q(\R[31][17] ), 
        .QN(n588) );
  DFFRX1 \R_reg[5][13]  ( .D(n2458), .CK(clk), .RN(reset_n), .Q(\R[5][13] ), 
        .QN(n1424) );
  DFFRX1 \R_reg[5][14]  ( .D(n2457), .CK(clk), .RN(reset_n), .Q(\R[5][14] ), 
        .QN(n1423) );
  DFFRX1 \R_reg[5][15]  ( .D(n2456), .CK(clk), .RN(reset_n), .Q(\R[5][15] ), 
        .QN(n1422) );
  DFFRX1 \R_reg[5][16]  ( .D(n2455), .CK(clk), .RN(reset_n), .Q(\R[5][16] ), 
        .QN(n1421) );
  DFFRX1 \R_reg[5][17]  ( .D(n2454), .CK(clk), .RN(reset_n), .Q(\R[5][17] ), 
        .QN(n1420) );
  DFFRX1 \R_reg[9][13]  ( .D(n2330), .CK(clk), .RN(reset_n), .Q(\R[9][13] ), 
        .QN(n1296) );
  DFFRX1 \R_reg[9][14]  ( .D(n2329), .CK(clk), .RN(reset_n), .Q(\R[9][14] ), 
        .QN(n1295) );
  DFFRX1 \R_reg[9][15]  ( .D(n2328), .CK(clk), .RN(reset_n), .Q(\R[9][15] ), 
        .QN(n1294) );
  DFFRX1 \R_reg[9][16]  ( .D(n2327), .CK(clk), .RN(reset_n), .Q(\R[9][16] ), 
        .QN(n1293) );
  DFFRX1 \R_reg[9][17]  ( .D(n2326), .CK(clk), .RN(reset_n), .Q(\R[9][17] ), 
        .QN(n1292) );
  DFFRX1 \R_reg[9][18]  ( .D(n2325), .CK(clk), .RN(reset_n), .Q(\R[9][18] ), 
        .QN(n1291) );
  DFFRX1 \R_reg[13][13]  ( .D(n2202), .CK(clk), .RN(reset_n), .Q(\R[13][13] ), 
        .QN(n1168) );
  DFFRX1 \R_reg[13][14]  ( .D(n2201), .CK(clk), .RN(reset_n), .Q(\R[13][14] ), 
        .QN(n1167) );
  DFFRX1 \R_reg[13][15]  ( .D(n2200), .CK(clk), .RN(reset_n), .Q(\R[13][15] ), 
        .QN(n1166) );
  DFFRX1 \R_reg[13][16]  ( .D(n2199), .CK(clk), .RN(reset_n), .Q(\R[13][16] ), 
        .QN(n1165) );
  DFFRX1 \R_reg[13][17]  ( .D(n2198), .CK(clk), .RN(reset_n), .Q(\R[13][17] ), 
        .QN(n1164) );
  DFFRX1 \R_reg[17][13]  ( .D(n2074), .CK(clk), .RN(reset_n), .Q(\R[17][13] ), 
        .QN(n1040) );
  DFFRX1 \R_reg[17][14]  ( .D(n2073), .CK(clk), .RN(reset_n), .Q(\R[17][14] ), 
        .QN(n1039) );
  DFFRX1 \R_reg[17][15]  ( .D(n2072), .CK(clk), .RN(reset_n), .Q(\R[17][15] ), 
        .QN(n1038) );
  DFFRX1 \R_reg[17][16]  ( .D(n2071), .CK(clk), .RN(reset_n), .Q(\R[17][16] ), 
        .QN(n1037) );
  DFFRX1 \R_reg[17][17]  ( .D(n2070), .CK(clk), .RN(reset_n), .Q(\R[17][17] ), 
        .QN(n1036) );
  DFFRX1 \R_reg[17][18]  ( .D(n2069), .CK(clk), .RN(reset_n), .Q(\R[17][18] ), 
        .QN(n1035) );
  DFFRX1 \R_reg[21][13]  ( .D(n1946), .CK(clk), .RN(reset_n), .Q(\R[21][13] ), 
        .QN(n912) );
  DFFRX1 \R_reg[21][14]  ( .D(n1945), .CK(clk), .RN(reset_n), .Q(\R[21][14] ), 
        .QN(n911) );
  DFFRX1 \R_reg[21][15]  ( .D(n1944), .CK(clk), .RN(reset_n), .Q(\R[21][15] ), 
        .QN(n910) );
  DFFRX1 \R_reg[21][16]  ( .D(n1943), .CK(clk), .RN(reset_n), .Q(\R[21][16] ), 
        .QN(n909) );
  DFFRX1 \R_reg[21][17]  ( .D(n1942), .CK(clk), .RN(reset_n), .Q(\R[21][17] ), 
        .QN(n908) );
  DFFRX1 \R_reg[25][13]  ( .D(n1818), .CK(clk), .RN(reset_n), .Q(\R[25][13] ), 
        .QN(n784) );
  DFFRX1 \R_reg[25][14]  ( .D(n1817), .CK(clk), .RN(reset_n), .Q(\R[25][14] ), 
        .QN(n783) );
  DFFRX1 \R_reg[25][15]  ( .D(n1816), .CK(clk), .RN(reset_n), .Q(\R[25][15] ), 
        .QN(n782) );
  DFFRX1 \R_reg[25][16]  ( .D(n1815), .CK(clk), .RN(reset_n), .Q(\R[25][16] ), 
        .QN(n781) );
  DFFRX1 \R_reg[25][17]  ( .D(n1814), .CK(clk), .RN(reset_n), .Q(\R[25][17] ), 
        .QN(n780) );
  DFFRX1 \R_reg[25][18]  ( .D(n1813), .CK(clk), .RN(reset_n), .Q(\R[25][18] ), 
        .QN(n779) );
  DFFRX1 \R_reg[29][13]  ( .D(n1690), .CK(clk), .RN(reset_n), .Q(\R[29][13] ), 
        .QN(n656) );
  DFFRX1 \R_reg[29][14]  ( .D(n1689), .CK(clk), .RN(reset_n), .Q(\R[29][14] ), 
        .QN(n655) );
  DFFRX1 \R_reg[29][15]  ( .D(n1688), .CK(clk), .RN(reset_n), .Q(\R[29][15] ), 
        .QN(n654) );
  DFFRX1 \R_reg[29][16]  ( .D(n1687), .CK(clk), .RN(reset_n), .Q(\R[29][16] ), 
        .QN(n653) );
  DFFRX1 \R_reg[29][17]  ( .D(n1686), .CK(clk), .RN(reset_n), .Q(\R[29][17] ), 
        .QN(n652) );
  DFFRX1 \R_reg[4][13]  ( .D(n2490), .CK(clk), .RN(reset_n), .Q(\R[4][13] ), 
        .QN(n1456) );
  DFFRX1 \R_reg[4][14]  ( .D(n2489), .CK(clk), .RN(reset_n), .Q(\R[4][14] ), 
        .QN(n1455) );
  DFFRX1 \R_reg[4][15]  ( .D(n2488), .CK(clk), .RN(reset_n), .Q(\R[4][15] ), 
        .QN(n1454) );
  DFFRX1 \R_reg[4][16]  ( .D(n2487), .CK(clk), .RN(reset_n), .Q(\R[4][16] ), 
        .QN(n1453) );
  DFFRX1 \R_reg[4][17]  ( .D(n2486), .CK(clk), .RN(reset_n), .Q(\R[4][17] ), 
        .QN(n1452) );
  DFFRX1 \R_reg[8][13]  ( .D(n2362), .CK(clk), .RN(reset_n), .Q(\R[8][13] ), 
        .QN(n1328) );
  DFFRX1 \R_reg[8][14]  ( .D(n2361), .CK(clk), .RN(reset_n), .Q(\R[8][14] ), 
        .QN(n1327) );
  DFFRX1 \R_reg[8][15]  ( .D(n2360), .CK(clk), .RN(reset_n), .Q(\R[8][15] ), 
        .QN(n1326) );
  DFFRX1 \R_reg[8][16]  ( .D(n2359), .CK(clk), .RN(reset_n), .Q(\R[8][16] ), 
        .QN(n1325) );
  DFFRX1 \R_reg[8][17]  ( .D(n2358), .CK(clk), .RN(reset_n), .Q(\R[8][17] ), 
        .QN(n1324) );
  DFFRX1 \R_reg[8][18]  ( .D(n2357), .CK(clk), .RN(reset_n), .Q(\R[8][18] ), 
        .QN(n1323) );
  DFFRX1 \R_reg[12][13]  ( .D(n2234), .CK(clk), .RN(reset_n), .Q(\R[12][13] ), 
        .QN(n1200) );
  DFFRX1 \R_reg[12][14]  ( .D(n2233), .CK(clk), .RN(reset_n), .Q(\R[12][14] ), 
        .QN(n1199) );
  DFFRX1 \R_reg[12][15]  ( .D(n2232), .CK(clk), .RN(reset_n), .Q(\R[12][15] ), 
        .QN(n1198) );
  DFFRX1 \R_reg[12][16]  ( .D(n2231), .CK(clk), .RN(reset_n), .Q(\R[12][16] ), 
        .QN(n1197) );
  DFFRX1 \R_reg[12][17]  ( .D(n2230), .CK(clk), .RN(reset_n), .Q(\R[12][17] ), 
        .QN(n1196) );
  DFFRX1 \R_reg[16][13]  ( .D(n2106), .CK(clk), .RN(reset_n), .Q(\R[16][13] ), 
        .QN(n1072) );
  DFFRX1 \R_reg[16][14]  ( .D(n2105), .CK(clk), .RN(reset_n), .Q(\R[16][14] ), 
        .QN(n1071) );
  DFFRX1 \R_reg[16][15]  ( .D(n2104), .CK(clk), .RN(reset_n), .Q(\R[16][15] ), 
        .QN(n1070) );
  DFFRX1 \R_reg[16][16]  ( .D(n2103), .CK(clk), .RN(reset_n), .Q(\R[16][16] ), 
        .QN(n1069) );
  DFFRX1 \R_reg[16][17]  ( .D(n2102), .CK(clk), .RN(reset_n), .Q(\R[16][17] ), 
        .QN(n1068) );
  DFFRX1 \R_reg[16][18]  ( .D(n2101), .CK(clk), .RN(reset_n), .Q(\R[16][18] ), 
        .QN(n1067) );
  DFFRX1 \R_reg[20][13]  ( .D(n1978), .CK(clk), .RN(reset_n), .Q(\R[20][13] ), 
        .QN(n944) );
  DFFRX1 \R_reg[20][14]  ( .D(n1977), .CK(clk), .RN(reset_n), .Q(\R[20][14] ), 
        .QN(n943) );
  DFFRX1 \R_reg[20][15]  ( .D(n1976), .CK(clk), .RN(reset_n), .Q(\R[20][15] ), 
        .QN(n942) );
  DFFRX1 \R_reg[20][16]  ( .D(n1975), .CK(clk), .RN(reset_n), .Q(\R[20][16] ), 
        .QN(n941) );
  DFFRX1 \R_reg[20][17]  ( .D(n1974), .CK(clk), .RN(reset_n), .Q(\R[20][17] ), 
        .QN(n940) );
  DFFRX1 \R_reg[24][13]  ( .D(n1850), .CK(clk), .RN(reset_n), .Q(\R[24][13] ), 
        .QN(n816) );
  DFFRX1 \R_reg[24][14]  ( .D(n1849), .CK(clk), .RN(reset_n), .Q(\R[24][14] ), 
        .QN(n815) );
  DFFRX1 \R_reg[24][15]  ( .D(n1848), .CK(clk), .RN(reset_n), .Q(\R[24][15] ), 
        .QN(n814) );
  DFFRX1 \R_reg[24][16]  ( .D(n1847), .CK(clk), .RN(reset_n), .Q(\R[24][16] ), 
        .QN(n813) );
  DFFRX1 \R_reg[24][17]  ( .D(n1846), .CK(clk), .RN(reset_n), .Q(\R[24][17] ), 
        .QN(n812) );
  DFFRX1 \R_reg[24][18]  ( .D(n1845), .CK(clk), .RN(reset_n), .Q(\R[24][18] ), 
        .QN(n811) );
  DFFRX1 \R_reg[28][13]  ( .D(n1722), .CK(clk), .RN(reset_n), .Q(\R[28][13] ), 
        .QN(n688) );
  DFFRX1 \R_reg[28][14]  ( .D(n1721), .CK(clk), .RN(reset_n), .Q(\R[28][14] ), 
        .QN(n687) );
  DFFRX1 \R_reg[28][15]  ( .D(n1720), .CK(clk), .RN(reset_n), .Q(\R[28][15] ), 
        .QN(n686) );
  DFFRX1 \R_reg[28][16]  ( .D(n1719), .CK(clk), .RN(reset_n), .Q(\R[28][16] ), 
        .QN(n685) );
  DFFRX1 \R_reg[28][17]  ( .D(n1718), .CK(clk), .RN(reset_n), .Q(\R[28][17] ), 
        .QN(n684) );
  DFFRX1 \R_reg[6][13]  ( .D(n2426), .CK(clk), .RN(reset_n), .Q(\R[6][13] ), 
        .QN(n1392) );
  DFFRX1 \R_reg[6][14]  ( .D(n2425), .CK(clk), .RN(reset_n), .Q(\R[6][14] ), 
        .QN(n1391) );
  DFFRX1 \R_reg[6][15]  ( .D(n2424), .CK(clk), .RN(reset_n), .Q(\R[6][15] ), 
        .QN(n1390) );
  DFFRX1 \R_reg[6][16]  ( .D(n2423), .CK(clk), .RN(reset_n), .Q(\R[6][16] ), 
        .QN(n1389) );
  DFFRX1 \R_reg[6][17]  ( .D(n2422), .CK(clk), .RN(reset_n), .Q(\R[6][17] ), 
        .QN(n1388) );
  DFFRX1 \R_reg[10][13]  ( .D(n2298), .CK(clk), .RN(reset_n), .Q(\R[10][13] ), 
        .QN(n1264) );
  DFFRX1 \R_reg[10][14]  ( .D(n2297), .CK(clk), .RN(reset_n), .Q(\R[10][14] ), 
        .QN(n1263) );
  DFFRX1 \R_reg[10][15]  ( .D(n2296), .CK(clk), .RN(reset_n), .Q(\R[10][15] ), 
        .QN(n1262) );
  DFFRX1 \R_reg[10][16]  ( .D(n2295), .CK(clk), .RN(reset_n), .Q(\R[10][16] ), 
        .QN(n1261) );
  DFFRX1 \R_reg[10][17]  ( .D(n2294), .CK(clk), .RN(reset_n), .Q(\R[10][17] ), 
        .QN(n1260) );
  DFFRX1 \R_reg[14][13]  ( .D(n2170), .CK(clk), .RN(reset_n), .Q(\R[14][13] ), 
        .QN(n1136) );
  DFFRX1 \R_reg[14][14]  ( .D(n2169), .CK(clk), .RN(reset_n), .Q(\R[14][14] ), 
        .QN(n1135) );
  DFFRX1 \R_reg[14][15]  ( .D(n2168), .CK(clk), .RN(reset_n), .Q(\R[14][15] ), 
        .QN(n1134) );
  DFFRX1 \R_reg[14][16]  ( .D(n2167), .CK(clk), .RN(reset_n), .Q(\R[14][16] ), 
        .QN(n1133) );
  DFFRX1 \R_reg[14][17]  ( .D(n2166), .CK(clk), .RN(reset_n), .Q(\R[14][17] ), 
        .QN(n1132) );
  DFFRX1 \R_reg[18][13]  ( .D(n2042), .CK(clk), .RN(reset_n), .Q(\R[18][13] ), 
        .QN(n1008) );
  DFFRX1 \R_reg[18][14]  ( .D(n2041), .CK(clk), .RN(reset_n), .Q(\R[18][14] ), 
        .QN(n1007) );
  DFFRX1 \R_reg[18][15]  ( .D(n2040), .CK(clk), .RN(reset_n), .Q(\R[18][15] ), 
        .QN(n1006) );
  DFFRX1 \R_reg[18][16]  ( .D(n2039), .CK(clk), .RN(reset_n), .Q(\R[18][16] ), 
        .QN(n1005) );
  DFFRX1 \R_reg[18][17]  ( .D(n2038), .CK(clk), .RN(reset_n), .Q(\R[18][17] ), 
        .QN(n1004) );
  DFFRX1 \R_reg[22][13]  ( .D(n1914), .CK(clk), .RN(reset_n), .Q(\R[22][13] ), 
        .QN(n880) );
  DFFRX1 \R_reg[22][14]  ( .D(n1913), .CK(clk), .RN(reset_n), .Q(\R[22][14] ), 
        .QN(n879) );
  DFFRX1 \R_reg[22][15]  ( .D(n1912), .CK(clk), .RN(reset_n), .Q(\R[22][15] ), 
        .QN(n878) );
  DFFRX1 \R_reg[22][16]  ( .D(n1911), .CK(clk), .RN(reset_n), .Q(\R[22][16] ), 
        .QN(n877) );
  DFFRX1 \R_reg[22][17]  ( .D(n1910), .CK(clk), .RN(reset_n), .Q(\R[22][17] ), 
        .QN(n876) );
  DFFRX1 \R_reg[26][13]  ( .D(n1786), .CK(clk), .RN(reset_n), .Q(\R[26][13] ), 
        .QN(n752) );
  DFFRX1 \R_reg[26][14]  ( .D(n1785), .CK(clk), .RN(reset_n), .Q(\R[26][14] ), 
        .QN(n751) );
  DFFRX1 \R_reg[26][15]  ( .D(n1784), .CK(clk), .RN(reset_n), .Q(\R[26][15] ), 
        .QN(n750) );
  DFFRX1 \R_reg[26][16]  ( .D(n1783), .CK(clk), .RN(reset_n), .Q(\R[26][16] ), 
        .QN(n749) );
  DFFRX1 \R_reg[26][17]  ( .D(n1782), .CK(clk), .RN(reset_n), .Q(\R[26][17] ), 
        .QN(n748) );
  DFFRX1 \R_reg[30][13]  ( .D(n1658), .CK(clk), .RN(reset_n), .Q(\R[30][13] ), 
        .QN(n624) );
  DFFRX1 \R_reg[30][14]  ( .D(n1657), .CK(clk), .RN(reset_n), .Q(\R[30][14] ), 
        .QN(n623) );
  DFFRX1 \R_reg[30][15]  ( .D(n1656), .CK(clk), .RN(reset_n), .Q(\R[30][15] ), 
        .QN(n622) );
  DFFRX1 \R_reg[30][16]  ( .D(n1655), .CK(clk), .RN(reset_n), .Q(\R[30][16] ), 
        .QN(n621) );
  DFFRX1 \R_reg[30][17]  ( .D(n1654), .CK(clk), .RN(reset_n), .Q(\R[30][17] ), 
        .QN(n620) );
  DFFRX1 \PC_reg[5]  ( .D(n2624), .CK(clk), .RN(reset_n), .Q(PC[5]), .QN(n1590) );
  DFFRX1 \PC_reg[6]  ( .D(n2623), .CK(clk), .RN(reset_n), .Q(PC[6]), .QN(n1589) );
  DFFRX1 \PC_reg[7]  ( .D(n2622), .CK(clk), .RN(reset_n), .Q(PC[7]), .QN(n1588) );
  DFFRX1 \PC_reg[8]  ( .D(n2621), .CK(clk), .RN(reset_n), .Q(PC[8]), .QN(n1587) );
  DFFRX1 \PC_reg[9]  ( .D(n2620), .CK(clk), .RN(reset_n), .Q(PC[9]), .QN(n1586) );
  DFFRX1 \PC_reg[10]  ( .D(n2619), .CK(clk), .RN(reset_n), .Q(PC[10]), .QN(
        n1585) );
  DFFRX1 \R_reg[1][12]  ( .D(n2587), .CK(clk), .RN(reset_n), .Q(\R[1][12] ), 
        .QN(n1553) );
  DFFRX1 \R_reg[1][13]  ( .D(n2586), .CK(clk), .RN(reset_n), .Q(\R[1][13] ), 
        .QN(n1552) );
  DFFRX1 \R_reg[1][14]  ( .D(n2585), .CK(clk), .RN(reset_n), .Q(\R[1][14] ), 
        .QN(n1551) );
  DFFRX1 \R_reg[1][15]  ( .D(n2584), .CK(clk), .RN(reset_n), .Q(\R[1][15] ), 
        .QN(n1550) );
  DFFRX1 \R_reg[1][16]  ( .D(n2583), .CK(clk), .RN(reset_n), .Q(\R[1][16] ), 
        .QN(n1549) );
  DFFRX1 \R_reg[1][17]  ( .D(n2582), .CK(clk), .RN(reset_n), .Q(\R[1][17] ), 
        .QN(n1548) );
  DFFRX1 \R_reg[3][13]  ( .D(n2522), .CK(clk), .RN(reset_n), .Q(\R[3][13] ), 
        .QN(n1488) );
  DFFRX1 \R_reg[3][14]  ( .D(n2521), .CK(clk), .RN(reset_n), .Q(\R[3][14] ), 
        .QN(n1487) );
  DFFRX1 \R_reg[3][15]  ( .D(n2520), .CK(clk), .RN(reset_n), .Q(\R[3][15] ), 
        .QN(n1486) );
  DFFRX1 \R_reg[3][16]  ( .D(n2519), .CK(clk), .RN(reset_n), .Q(\R[3][16] ), 
        .QN(n1485) );
  DFFRX1 \R_reg[3][17]  ( .D(n2518), .CK(clk), .RN(reset_n), .Q(\R[3][17] ), 
        .QN(n1484) );
  DFFRX1 \R_reg[2][13]  ( .D(n2554), .CK(clk), .RN(reset_n), .QN(n1520) );
  DFFRX1 \R_reg[2][14]  ( .D(n2553), .CK(clk), .RN(reset_n), .QN(n1519) );
  DFFRX1 \R_reg[2][15]  ( .D(n2552), .CK(clk), .RN(reset_n), .QN(n1518) );
  DFFRX1 \R_reg[2][16]  ( .D(n2551), .CK(clk), .RN(reset_n), .QN(n1517) );
  DFFRX1 \R_reg[2][17]  ( .D(n2550), .CK(clk), .RN(reset_n), .QN(n1516) );
  DFFRX1 \counter_reg[1]  ( .D(N127), .CK(clk), .RN(reset_n), .Q(counter[1])
         );
  DFFRX1 \counter_reg[0]  ( .D(N126), .CK(clk), .RN(reset_n), .Q(counter[0])
         );
  DFFRX1 \R_reg[7][7]  ( .D(n2400), .CK(clk), .RN(reset_n), .Q(\R[7][7] ), 
        .QN(n1366) );
  DFFRX1 \R_reg[7][8]  ( .D(n2399), .CK(clk), .RN(reset_n), .Q(\R[7][8] ), 
        .QN(n1365) );
  DFFRX1 \R_reg[7][9]  ( .D(n2398), .CK(clk), .RN(reset_n), .Q(\R[7][9] ), 
        .QN(n1364) );
  DFFRX1 \R_reg[7][10]  ( .D(n2397), .CK(clk), .RN(reset_n), .Q(\R[7][10] ), 
        .QN(n1363) );
  DFFRX1 \R_reg[7][11]  ( .D(n2396), .CK(clk), .RN(reset_n), .Q(\R[7][11] ), 
        .QN(n1362) );
  DFFRX1 \R_reg[7][12]  ( .D(n2395), .CK(clk), .RN(reset_n), .Q(\R[7][12] ), 
        .QN(n1361) );
  DFFRX1 \R_reg[11][7]  ( .D(n2272), .CK(clk), .RN(reset_n), .Q(\R[11][7] ), 
        .QN(n1238) );
  DFFRX1 \R_reg[11][8]  ( .D(n2271), .CK(clk), .RN(reset_n), .Q(\R[11][8] ), 
        .QN(n1237) );
  DFFRX1 \R_reg[11][9]  ( .D(n2270), .CK(clk), .RN(reset_n), .Q(\R[11][9] ), 
        .QN(n1236) );
  DFFRX1 \R_reg[11][10]  ( .D(n2269), .CK(clk), .RN(reset_n), .Q(\R[11][10] ), 
        .QN(n1235) );
  DFFRX1 \R_reg[11][11]  ( .D(n2268), .CK(clk), .RN(reset_n), .Q(\R[11][11] ), 
        .QN(n1234) );
  DFFRX1 \R_reg[11][12]  ( .D(n2267), .CK(clk), .RN(reset_n), .Q(\R[11][12] ), 
        .QN(n1233) );
  DFFRX1 \R_reg[15][7]  ( .D(n2144), .CK(clk), .RN(reset_n), .Q(\R[15][7] ), 
        .QN(n1110) );
  DFFRX1 \R_reg[15][8]  ( .D(n2143), .CK(clk), .RN(reset_n), .Q(\R[15][8] ), 
        .QN(n1109) );
  DFFRX1 \R_reg[15][9]  ( .D(n2142), .CK(clk), .RN(reset_n), .Q(\R[15][9] ), 
        .QN(n1108) );
  DFFRX1 \R_reg[15][10]  ( .D(n2141), .CK(clk), .RN(reset_n), .Q(\R[15][10] ), 
        .QN(n1107) );
  DFFRX1 \R_reg[15][11]  ( .D(n2140), .CK(clk), .RN(reset_n), .Q(\R[15][11] ), 
        .QN(n1106) );
  DFFRX1 \R_reg[15][12]  ( .D(n2139), .CK(clk), .RN(reset_n), .Q(\R[15][12] ), 
        .QN(n1105) );
  DFFRX1 \R_reg[19][7]  ( .D(n2016), .CK(clk), .RN(reset_n), .Q(\R[19][7] ), 
        .QN(n982) );
  DFFRX1 \R_reg[19][8]  ( .D(n2015), .CK(clk), .RN(reset_n), .Q(\R[19][8] ), 
        .QN(n981) );
  DFFRX1 \R_reg[19][9]  ( .D(n2014), .CK(clk), .RN(reset_n), .Q(\R[19][9] ), 
        .QN(n980) );
  DFFRX1 \R_reg[19][10]  ( .D(n2013), .CK(clk), .RN(reset_n), .Q(\R[19][10] ), 
        .QN(n979) );
  DFFRX1 \R_reg[19][11]  ( .D(n2012), .CK(clk), .RN(reset_n), .Q(\R[19][11] ), 
        .QN(n978) );
  DFFRX1 \R_reg[19][12]  ( .D(n2011), .CK(clk), .RN(reset_n), .Q(\R[19][12] ), 
        .QN(n977) );
  DFFRX1 \R_reg[23][7]  ( .D(n1888), .CK(clk), .RN(reset_n), .Q(\R[23][7] ), 
        .QN(n854) );
  DFFRX1 \R_reg[23][8]  ( .D(n1887), .CK(clk), .RN(reset_n), .Q(\R[23][8] ), 
        .QN(n853) );
  DFFRX1 \R_reg[23][9]  ( .D(n1886), .CK(clk), .RN(reset_n), .Q(\R[23][9] ), 
        .QN(n852) );
  DFFRX1 \R_reg[23][10]  ( .D(n1885), .CK(clk), .RN(reset_n), .Q(\R[23][10] ), 
        .QN(n851) );
  DFFRX1 \R_reg[23][11]  ( .D(n1884), .CK(clk), .RN(reset_n), .Q(\R[23][11] ), 
        .QN(n850) );
  DFFRX1 \R_reg[23][12]  ( .D(n1883), .CK(clk), .RN(reset_n), .Q(\R[23][12] ), 
        .QN(n849) );
  DFFRX1 \R_reg[27][7]  ( .D(n1760), .CK(clk), .RN(reset_n), .Q(\R[27][7] ), 
        .QN(n726) );
  DFFRX1 \R_reg[27][8]  ( .D(n1759), .CK(clk), .RN(reset_n), .Q(\R[27][8] ), 
        .QN(n725) );
  DFFRX1 \R_reg[27][9]  ( .D(n1758), .CK(clk), .RN(reset_n), .Q(\R[27][9] ), 
        .QN(n724) );
  DFFRX1 \R_reg[27][10]  ( .D(n1757), .CK(clk), .RN(reset_n), .Q(\R[27][10] ), 
        .QN(n723) );
  DFFRX1 \R_reg[27][11]  ( .D(n1756), .CK(clk), .RN(reset_n), .Q(\R[27][11] ), 
        .QN(n722) );
  DFFRX1 \R_reg[27][12]  ( .D(n1755), .CK(clk), .RN(reset_n), .Q(\R[27][12] ), 
        .QN(n721) );
  DFFRX1 \R_reg[31][7]  ( .D(n1632), .CK(clk), .RN(reset_n), .Q(\R[31][7] ), 
        .QN(n598) );
  DFFRX1 \R_reg[31][8]  ( .D(n1631), .CK(clk), .RN(reset_n), .Q(\R[31][8] ), 
        .QN(n597) );
  DFFRX1 \R_reg[31][9]  ( .D(n1630), .CK(clk), .RN(reset_n), .Q(\R[31][9] ), 
        .QN(n596) );
  DFFRX1 \R_reg[31][10]  ( .D(n1629), .CK(clk), .RN(reset_n), .Q(\R[31][10] ), 
        .QN(n595) );
  DFFRX1 \R_reg[31][11]  ( .D(n1628), .CK(clk), .RN(reset_n), .Q(\R[31][11] ), 
        .QN(n594) );
  DFFRX1 \R_reg[31][12]  ( .D(n1627), .CK(clk), .RN(reset_n), .Q(\R[31][12] ), 
        .QN(n593) );
  DFFRX1 \R_reg[5][7]  ( .D(n2464), .CK(clk), .RN(reset_n), .Q(\R[5][7] ), 
        .QN(n1430) );
  DFFRX1 \R_reg[5][8]  ( .D(n2463), .CK(clk), .RN(reset_n), .Q(\R[5][8] ), 
        .QN(n1429) );
  DFFRX1 \R_reg[5][9]  ( .D(n2462), .CK(clk), .RN(reset_n), .Q(\R[5][9] ), 
        .QN(n1428) );
  DFFRX1 \R_reg[5][10]  ( .D(n2461), .CK(clk), .RN(reset_n), .Q(\R[5][10] ), 
        .QN(n1427) );
  DFFRX1 \R_reg[5][11]  ( .D(n2460), .CK(clk), .RN(reset_n), .Q(\R[5][11] ), 
        .QN(n1426) );
  DFFRX1 \R_reg[5][12]  ( .D(n2459), .CK(clk), .RN(reset_n), .Q(\R[5][12] ), 
        .QN(n1425) );
  DFFRX1 \R_reg[9][7]  ( .D(n2336), .CK(clk), .RN(reset_n), .Q(\R[9][7] ), 
        .QN(n1302) );
  DFFRX1 \R_reg[9][8]  ( .D(n2335), .CK(clk), .RN(reset_n), .Q(\R[9][8] ), 
        .QN(n1301) );
  DFFRX1 \R_reg[9][9]  ( .D(n2334), .CK(clk), .RN(reset_n), .Q(\R[9][9] ), 
        .QN(n1300) );
  DFFRX1 \R_reg[9][10]  ( .D(n2333), .CK(clk), .RN(reset_n), .Q(\R[9][10] ), 
        .QN(n1299) );
  DFFRX1 \R_reg[9][11]  ( .D(n2332), .CK(clk), .RN(reset_n), .Q(\R[9][11] ), 
        .QN(n1298) );
  DFFRX1 \R_reg[9][12]  ( .D(n2331), .CK(clk), .RN(reset_n), .Q(\R[9][12] ), 
        .QN(n1297) );
  DFFRX1 \R_reg[13][7]  ( .D(n2208), .CK(clk), .RN(reset_n), .Q(\R[13][7] ), 
        .QN(n1174) );
  DFFRX1 \R_reg[13][8]  ( .D(n2207), .CK(clk), .RN(reset_n), .Q(\R[13][8] ), 
        .QN(n1173) );
  DFFRX1 \R_reg[13][9]  ( .D(n2206), .CK(clk), .RN(reset_n), .Q(\R[13][9] ), 
        .QN(n1172) );
  DFFRX1 \R_reg[13][10]  ( .D(n2205), .CK(clk), .RN(reset_n), .Q(\R[13][10] ), 
        .QN(n1171) );
  DFFRX1 \R_reg[13][11]  ( .D(n2204), .CK(clk), .RN(reset_n), .Q(\R[13][11] ), 
        .QN(n1170) );
  DFFRX1 \R_reg[13][12]  ( .D(n2203), .CK(clk), .RN(reset_n), .Q(\R[13][12] ), 
        .QN(n1169) );
  DFFRX1 \R_reg[17][7]  ( .D(n2080), .CK(clk), .RN(reset_n), .Q(\R[17][7] ), 
        .QN(n1046) );
  DFFRX1 \R_reg[17][8]  ( .D(n2079), .CK(clk), .RN(reset_n), .Q(\R[17][8] ), 
        .QN(n1045) );
  DFFRX1 \R_reg[17][9]  ( .D(n2078), .CK(clk), .RN(reset_n), .Q(\R[17][9] ), 
        .QN(n1044) );
  DFFRX1 \R_reg[17][10]  ( .D(n2077), .CK(clk), .RN(reset_n), .Q(\R[17][10] ), 
        .QN(n1043) );
  DFFRX1 \R_reg[17][11]  ( .D(n2076), .CK(clk), .RN(reset_n), .Q(\R[17][11] ), 
        .QN(n1042) );
  DFFRX1 \R_reg[17][12]  ( .D(n2075), .CK(clk), .RN(reset_n), .Q(\R[17][12] ), 
        .QN(n1041) );
  DFFRX1 \R_reg[21][7]  ( .D(n1952), .CK(clk), .RN(reset_n), .Q(\R[21][7] ), 
        .QN(n918) );
  DFFRX1 \R_reg[21][8]  ( .D(n1951), .CK(clk), .RN(reset_n), .Q(\R[21][8] ), 
        .QN(n917) );
  DFFRX1 \R_reg[21][9]  ( .D(n1950), .CK(clk), .RN(reset_n), .Q(\R[21][9] ), 
        .QN(n916) );
  DFFRX1 \R_reg[21][10]  ( .D(n1949), .CK(clk), .RN(reset_n), .Q(\R[21][10] ), 
        .QN(n915) );
  DFFRX1 \R_reg[21][11]  ( .D(n1948), .CK(clk), .RN(reset_n), .Q(\R[21][11] ), 
        .QN(n914) );
  DFFRX1 \R_reg[21][12]  ( .D(n1947), .CK(clk), .RN(reset_n), .Q(\R[21][12] ), 
        .QN(n913) );
  DFFRX1 \R_reg[25][7]  ( .D(n1824), .CK(clk), .RN(reset_n), .Q(\R[25][7] ), 
        .QN(n790) );
  DFFRX1 \R_reg[25][8]  ( .D(n1823), .CK(clk), .RN(reset_n), .Q(\R[25][8] ), 
        .QN(n789) );
  DFFRX1 \R_reg[25][9]  ( .D(n1822), .CK(clk), .RN(reset_n), .Q(\R[25][9] ), 
        .QN(n788) );
  DFFRX1 \R_reg[25][10]  ( .D(n1821), .CK(clk), .RN(reset_n), .Q(\R[25][10] ), 
        .QN(n787) );
  DFFRX1 \R_reg[25][11]  ( .D(n1820), .CK(clk), .RN(reset_n), .Q(\R[25][11] ), 
        .QN(n786) );
  DFFRX1 \R_reg[25][12]  ( .D(n1819), .CK(clk), .RN(reset_n), .Q(\R[25][12] ), 
        .QN(n785) );
  DFFRX1 \R_reg[29][7]  ( .D(n1696), .CK(clk), .RN(reset_n), .Q(\R[29][7] ), 
        .QN(n662) );
  DFFRX1 \R_reg[29][8]  ( .D(n1695), .CK(clk), .RN(reset_n), .Q(\R[29][8] ), 
        .QN(n661) );
  DFFRX1 \R_reg[29][9]  ( .D(n1694), .CK(clk), .RN(reset_n), .Q(\R[29][9] ), 
        .QN(n660) );
  DFFRX1 \R_reg[29][10]  ( .D(n1693), .CK(clk), .RN(reset_n), .Q(\R[29][10] ), 
        .QN(n659) );
  DFFRX1 \R_reg[29][11]  ( .D(n1692), .CK(clk), .RN(reset_n), .Q(\R[29][11] ), 
        .QN(n658) );
  DFFRX1 \R_reg[29][12]  ( .D(n1691), .CK(clk), .RN(reset_n), .Q(\R[29][12] ), 
        .QN(n657) );
  DFFRX1 \R_reg[4][7]  ( .D(n2496), .CK(clk), .RN(reset_n), .Q(\R[4][7] ), 
        .QN(n1462) );
  DFFRX1 \R_reg[4][8]  ( .D(n2495), .CK(clk), .RN(reset_n), .Q(\R[4][8] ), 
        .QN(n1461) );
  DFFRX1 \R_reg[4][9]  ( .D(n2494), .CK(clk), .RN(reset_n), .Q(\R[4][9] ), 
        .QN(n1460) );
  DFFRX1 \R_reg[4][10]  ( .D(n2493), .CK(clk), .RN(reset_n), .Q(\R[4][10] ), 
        .QN(n1459) );
  DFFRX1 \R_reg[4][11]  ( .D(n2492), .CK(clk), .RN(reset_n), .Q(\R[4][11] ), 
        .QN(n1458) );
  DFFRX1 \R_reg[4][12]  ( .D(n2491), .CK(clk), .RN(reset_n), .Q(\R[4][12] ), 
        .QN(n1457) );
  DFFRX1 \R_reg[8][7]  ( .D(n2368), .CK(clk), .RN(reset_n), .Q(\R[8][7] ), 
        .QN(n1334) );
  DFFRX1 \R_reg[8][8]  ( .D(n2367), .CK(clk), .RN(reset_n), .Q(\R[8][8] ), 
        .QN(n1333) );
  DFFRX1 \R_reg[8][9]  ( .D(n2366), .CK(clk), .RN(reset_n), .Q(\R[8][9] ), 
        .QN(n1332) );
  DFFRX1 \R_reg[8][10]  ( .D(n2365), .CK(clk), .RN(reset_n), .Q(\R[8][10] ), 
        .QN(n1331) );
  DFFRX1 \R_reg[8][11]  ( .D(n2364), .CK(clk), .RN(reset_n), .Q(\R[8][11] ), 
        .QN(n1330) );
  DFFRX1 \R_reg[8][12]  ( .D(n2363), .CK(clk), .RN(reset_n), .Q(\R[8][12] ), 
        .QN(n1329) );
  DFFRX1 \R_reg[12][7]  ( .D(n2240), .CK(clk), .RN(reset_n), .Q(\R[12][7] ), 
        .QN(n1206) );
  DFFRX1 \R_reg[12][8]  ( .D(n2239), .CK(clk), .RN(reset_n), .Q(\R[12][8] ), 
        .QN(n1205) );
  DFFRX1 \R_reg[12][9]  ( .D(n2238), .CK(clk), .RN(reset_n), .Q(\R[12][9] ), 
        .QN(n1204) );
  DFFRX1 \R_reg[12][10]  ( .D(n2237), .CK(clk), .RN(reset_n), .Q(\R[12][10] ), 
        .QN(n1203) );
  DFFRX1 \R_reg[12][11]  ( .D(n2236), .CK(clk), .RN(reset_n), .Q(\R[12][11] ), 
        .QN(n1202) );
  DFFRX1 \R_reg[12][12]  ( .D(n2235), .CK(clk), .RN(reset_n), .Q(\R[12][12] ), 
        .QN(n1201) );
  DFFRX1 \R_reg[16][7]  ( .D(n2112), .CK(clk), .RN(reset_n), .Q(\R[16][7] ), 
        .QN(n1078) );
  DFFRX1 \R_reg[16][8]  ( .D(n2111), .CK(clk), .RN(reset_n), .Q(\R[16][8] ), 
        .QN(n1077) );
  DFFRX1 \R_reg[16][9]  ( .D(n2110), .CK(clk), .RN(reset_n), .Q(\R[16][9] ), 
        .QN(n1076) );
  DFFRX1 \R_reg[16][10]  ( .D(n2109), .CK(clk), .RN(reset_n), .Q(\R[16][10] ), 
        .QN(n1075) );
  DFFRX1 \R_reg[16][11]  ( .D(n2108), .CK(clk), .RN(reset_n), .Q(\R[16][11] ), 
        .QN(n1074) );
  DFFRX1 \R_reg[16][12]  ( .D(n2107), .CK(clk), .RN(reset_n), .Q(\R[16][12] ), 
        .QN(n1073) );
  DFFRX1 \R_reg[20][7]  ( .D(n1984), .CK(clk), .RN(reset_n), .Q(\R[20][7] ), 
        .QN(n950) );
  DFFRX1 \R_reg[20][8]  ( .D(n1983), .CK(clk), .RN(reset_n), .Q(\R[20][8] ), 
        .QN(n949) );
  DFFRX1 \R_reg[20][9]  ( .D(n1982), .CK(clk), .RN(reset_n), .Q(\R[20][9] ), 
        .QN(n948) );
  DFFRX1 \R_reg[20][10]  ( .D(n1981), .CK(clk), .RN(reset_n), .Q(\R[20][10] ), 
        .QN(n947) );
  DFFRX1 \R_reg[20][11]  ( .D(n1980), .CK(clk), .RN(reset_n), .Q(\R[20][11] ), 
        .QN(n946) );
  DFFRX1 \R_reg[20][12]  ( .D(n1979), .CK(clk), .RN(reset_n), .Q(\R[20][12] ), 
        .QN(n945) );
  DFFRX1 \R_reg[24][7]  ( .D(n1856), .CK(clk), .RN(reset_n), .Q(\R[24][7] ), 
        .QN(n822) );
  DFFRX1 \R_reg[24][8]  ( .D(n1855), .CK(clk), .RN(reset_n), .Q(\R[24][8] ), 
        .QN(n821) );
  DFFRX1 \R_reg[24][9]  ( .D(n1854), .CK(clk), .RN(reset_n), .Q(\R[24][9] ), 
        .QN(n820) );
  DFFRX1 \R_reg[24][10]  ( .D(n1853), .CK(clk), .RN(reset_n), .Q(\R[24][10] ), 
        .QN(n819) );
  DFFRX1 \R_reg[24][11]  ( .D(n1852), .CK(clk), .RN(reset_n), .Q(\R[24][11] ), 
        .QN(n818) );
  DFFRX1 \R_reg[24][12]  ( .D(n1851), .CK(clk), .RN(reset_n), .Q(\R[24][12] ), 
        .QN(n817) );
  DFFRX1 \R_reg[28][7]  ( .D(n1728), .CK(clk), .RN(reset_n), .Q(\R[28][7] ), 
        .QN(n694) );
  DFFRX1 \R_reg[28][8]  ( .D(n1727), .CK(clk), .RN(reset_n), .Q(\R[28][8] ), 
        .QN(n693) );
  DFFRX1 \R_reg[28][9]  ( .D(n1726), .CK(clk), .RN(reset_n), .Q(\R[28][9] ), 
        .QN(n692) );
  DFFRX1 \R_reg[28][10]  ( .D(n1725), .CK(clk), .RN(reset_n), .Q(\R[28][10] ), 
        .QN(n691) );
  DFFRX1 \R_reg[28][11]  ( .D(n1724), .CK(clk), .RN(reset_n), .Q(\R[28][11] ), 
        .QN(n690) );
  DFFRX1 \R_reg[28][12]  ( .D(n1723), .CK(clk), .RN(reset_n), .Q(\R[28][12] ), 
        .QN(n689) );
  DFFRX1 \R_reg[6][7]  ( .D(n2432), .CK(clk), .RN(reset_n), .Q(\R[6][7] ), 
        .QN(n1398) );
  DFFRX1 \R_reg[6][8]  ( .D(n2431), .CK(clk), .RN(reset_n), .Q(\R[6][8] ), 
        .QN(n1397) );
  DFFRX1 \R_reg[6][9]  ( .D(n2430), .CK(clk), .RN(reset_n), .Q(\R[6][9] ), 
        .QN(n1396) );
  DFFRX1 \R_reg[6][10]  ( .D(n2429), .CK(clk), .RN(reset_n), .Q(\R[6][10] ), 
        .QN(n1395) );
  DFFRX1 \R_reg[6][11]  ( .D(n2428), .CK(clk), .RN(reset_n), .Q(\R[6][11] ), 
        .QN(n1394) );
  DFFRX1 \R_reg[6][12]  ( .D(n2427), .CK(clk), .RN(reset_n), .Q(\R[6][12] ), 
        .QN(n1393) );
  DFFRX1 \R_reg[10][7]  ( .D(n2304), .CK(clk), .RN(reset_n), .Q(\R[10][7] ), 
        .QN(n1270) );
  DFFRX1 \R_reg[10][8]  ( .D(n2303), .CK(clk), .RN(reset_n), .Q(\R[10][8] ), 
        .QN(n1269) );
  DFFRX1 \R_reg[10][9]  ( .D(n2302), .CK(clk), .RN(reset_n), .Q(\R[10][9] ), 
        .QN(n1268) );
  DFFRX1 \R_reg[10][10]  ( .D(n2301), .CK(clk), .RN(reset_n), .Q(\R[10][10] ), 
        .QN(n1267) );
  DFFRX1 \R_reg[10][11]  ( .D(n2300), .CK(clk), .RN(reset_n), .Q(\R[10][11] ), 
        .QN(n1266) );
  DFFRX1 \R_reg[10][12]  ( .D(n2299), .CK(clk), .RN(reset_n), .Q(\R[10][12] ), 
        .QN(n1265) );
  DFFRX1 \R_reg[14][7]  ( .D(n2176), .CK(clk), .RN(reset_n), .Q(\R[14][7] ), 
        .QN(n1142) );
  DFFRX1 \R_reg[14][8]  ( .D(n2175), .CK(clk), .RN(reset_n), .Q(\R[14][8] ), 
        .QN(n1141) );
  DFFRX1 \R_reg[14][9]  ( .D(n2174), .CK(clk), .RN(reset_n), .Q(\R[14][9] ), 
        .QN(n1140) );
  DFFRX1 \R_reg[14][10]  ( .D(n2173), .CK(clk), .RN(reset_n), .Q(\R[14][10] ), 
        .QN(n1139) );
  DFFRX1 \R_reg[14][11]  ( .D(n2172), .CK(clk), .RN(reset_n), .Q(\R[14][11] ), 
        .QN(n1138) );
  DFFRX1 \R_reg[14][12]  ( .D(n2171), .CK(clk), .RN(reset_n), .Q(\R[14][12] ), 
        .QN(n1137) );
  DFFRX1 \R_reg[18][7]  ( .D(n2048), .CK(clk), .RN(reset_n), .Q(\R[18][7] ), 
        .QN(n1014) );
  DFFRX1 \R_reg[18][8]  ( .D(n2047), .CK(clk), .RN(reset_n), .Q(\R[18][8] ), 
        .QN(n1013) );
  DFFRX1 \R_reg[18][9]  ( .D(n2046), .CK(clk), .RN(reset_n), .Q(\R[18][9] ), 
        .QN(n1012) );
  DFFRX1 \R_reg[18][10]  ( .D(n2045), .CK(clk), .RN(reset_n), .Q(\R[18][10] ), 
        .QN(n1011) );
  DFFRX1 \R_reg[18][11]  ( .D(n2044), .CK(clk), .RN(reset_n), .Q(\R[18][11] ), 
        .QN(n1010) );
  DFFRX1 \R_reg[18][12]  ( .D(n2043), .CK(clk), .RN(reset_n), .Q(\R[18][12] ), 
        .QN(n1009) );
  DFFRX1 \R_reg[22][7]  ( .D(n1920), .CK(clk), .RN(reset_n), .Q(\R[22][7] ), 
        .QN(n886) );
  DFFRX1 \R_reg[22][8]  ( .D(n1919), .CK(clk), .RN(reset_n), .Q(\R[22][8] ), 
        .QN(n885) );
  DFFRX1 \R_reg[22][9]  ( .D(n1918), .CK(clk), .RN(reset_n), .Q(\R[22][9] ), 
        .QN(n884) );
  DFFRX1 \R_reg[22][10]  ( .D(n1917), .CK(clk), .RN(reset_n), .Q(\R[22][10] ), 
        .QN(n883) );
  DFFRX1 \R_reg[22][11]  ( .D(n1916), .CK(clk), .RN(reset_n), .Q(\R[22][11] ), 
        .QN(n882) );
  DFFRX1 \R_reg[22][12]  ( .D(n1915), .CK(clk), .RN(reset_n), .Q(\R[22][12] ), 
        .QN(n881) );
  DFFRX1 \R_reg[26][7]  ( .D(n1792), .CK(clk), .RN(reset_n), .Q(\R[26][7] ), 
        .QN(n758) );
  DFFRX1 \R_reg[26][8]  ( .D(n1791), .CK(clk), .RN(reset_n), .Q(\R[26][8] ), 
        .QN(n757) );
  DFFRX1 \R_reg[26][9]  ( .D(n1790), .CK(clk), .RN(reset_n), .Q(\R[26][9] ), 
        .QN(n756) );
  DFFRX1 \R_reg[26][10]  ( .D(n1789), .CK(clk), .RN(reset_n), .Q(\R[26][10] ), 
        .QN(n755) );
  DFFRX1 \R_reg[26][11]  ( .D(n1788), .CK(clk), .RN(reset_n), .Q(\R[26][11] ), 
        .QN(n754) );
  DFFRX1 \R_reg[26][12]  ( .D(n1787), .CK(clk), .RN(reset_n), .Q(\R[26][12] ), 
        .QN(n753) );
  DFFRX1 \R_reg[30][7]  ( .D(n1664), .CK(clk), .RN(reset_n), .Q(\R[30][7] ), 
        .QN(n630) );
  DFFRX1 \R_reg[30][8]  ( .D(n1663), .CK(clk), .RN(reset_n), .Q(\R[30][8] ), 
        .QN(n629) );
  DFFRX1 \R_reg[30][9]  ( .D(n1662), .CK(clk), .RN(reset_n), .Q(\R[30][9] ), 
        .QN(n628) );
  DFFRX1 \R_reg[30][10]  ( .D(n1661), .CK(clk), .RN(reset_n), .Q(\R[30][10] ), 
        .QN(n627) );
  DFFRX1 \R_reg[30][11]  ( .D(n1660), .CK(clk), .RN(reset_n), .Q(\R[30][11] ), 
        .QN(n626) );
  DFFRX1 \R_reg[30][12]  ( .D(n1659), .CK(clk), .RN(reset_n), .Q(\R[30][12] ), 
        .QN(n625) );
  DFFRX1 \PC_reg[1]  ( .D(n2628), .CK(clk), .RN(reset_n), .Q(PC[1]), .QN(n1594) );
  DFFRX1 \PC_reg[2]  ( .D(n2627), .CK(clk), .RN(reset_n), .Q(PC[2]), .QN(n1593) );
  DFFRX1 \PC_reg[3]  ( .D(n2626), .CK(clk), .RN(reset_n), .Q(PC[3]), .QN(n1592) );
  DFFRX1 \PC_reg[4]  ( .D(n2625), .CK(clk), .RN(reset_n), .Q(PC[4]), .QN(n1591) );
  DFFRX1 \R_reg[1][7]  ( .D(n2592), .CK(clk), .RN(reset_n), .Q(\R[1][7] ), 
        .QN(n1558) );
  DFFRX1 \R_reg[1][8]  ( .D(n2591), .CK(clk), .RN(reset_n), .Q(\R[1][8] ), 
        .QN(n1557) );
  DFFRX1 \R_reg[1][9]  ( .D(n2590), .CK(clk), .RN(reset_n), .Q(\R[1][9] ), 
        .QN(n1556) );
  DFFRX1 \R_reg[1][10]  ( .D(n2589), .CK(clk), .RN(reset_n), .Q(\R[1][10] ), 
        .QN(n1555) );
  DFFRX1 \R_reg[1][11]  ( .D(n2588), .CK(clk), .RN(reset_n), .Q(\R[1][11] ), 
        .QN(n1554) );
  DFFRX1 \R_reg[3][7]  ( .D(n2528), .CK(clk), .RN(reset_n), .Q(\R[3][7] ), 
        .QN(n1494) );
  DFFRX1 \R_reg[3][8]  ( .D(n2527), .CK(clk), .RN(reset_n), .Q(\R[3][8] ), 
        .QN(n1493) );
  DFFRX1 \R_reg[3][9]  ( .D(n2526), .CK(clk), .RN(reset_n), .Q(\R[3][9] ), 
        .QN(n1492) );
  DFFRX1 \R_reg[3][10]  ( .D(n2525), .CK(clk), .RN(reset_n), .Q(\R[3][10] ), 
        .QN(n1491) );
  DFFRX1 \R_reg[3][11]  ( .D(n2524), .CK(clk), .RN(reset_n), .Q(\R[3][11] ), 
        .QN(n1490) );
  DFFRX1 \R_reg[3][12]  ( .D(n2523), .CK(clk), .RN(reset_n), .Q(\R[3][12] ), 
        .QN(n1489) );
  DFFRX1 \R_reg[2][7]  ( .D(n2560), .CK(clk), .RN(reset_n), .QN(n1526) );
  DFFRX1 \R_reg[2][8]  ( .D(n2559), .CK(clk), .RN(reset_n), .QN(n1525) );
  DFFRX1 \R_reg[2][9]  ( .D(n2558), .CK(clk), .RN(reset_n), .QN(n1524) );
  DFFRX1 \R_reg[2][10]  ( .D(n2557), .CK(clk), .RN(reset_n), .QN(n1523) );
  DFFRX1 \R_reg[2][11]  ( .D(n2556), .CK(clk), .RN(reset_n), .QN(n1522) );
  DFFRX1 \R_reg[2][12]  ( .D(n2555), .CK(clk), .RN(reset_n), .QN(n1521) );
  DFFRX1 \PC_reg[0]  ( .D(n2629), .CK(clk), .RN(reset_n), .Q(PC[0]), .QN(n1595) );
  DFFRX1 \R_reg[7][0]  ( .D(n2407), .CK(clk), .RN(reset_n), .Q(\R[7][0] ), 
        .QN(n1373) );
  DFFRX1 \R_reg[7][1]  ( .D(n2406), .CK(clk), .RN(reset_n), .Q(\R[7][1] ), 
        .QN(n1372) );
  DFFRX1 \R_reg[7][2]  ( .D(n2405), .CK(clk), .RN(reset_n), .Q(\R[7][2] ), 
        .QN(n1371) );
  DFFRX1 \R_reg[7][3]  ( .D(n2404), .CK(clk), .RN(reset_n), .Q(\R[7][3] ), 
        .QN(n1370) );
  DFFRX1 \R_reg[7][4]  ( .D(n2403), .CK(clk), .RN(reset_n), .Q(\R[7][4] ), 
        .QN(n1369) );
  DFFRX1 \R_reg[7][5]  ( .D(n2402), .CK(clk), .RN(reset_n), .Q(\R[7][5] ), 
        .QN(n1368) );
  DFFRX1 \R_reg[7][6]  ( .D(n2401), .CK(clk), .RN(reset_n), .Q(\R[7][6] ), 
        .QN(n1367) );
  DFFRX1 \R_reg[11][0]  ( .D(n2279), .CK(clk), .RN(reset_n), .Q(\R[11][0] ), 
        .QN(n1245) );
  DFFRX1 \R_reg[11][1]  ( .D(n2278), .CK(clk), .RN(reset_n), .Q(\R[11][1] ), 
        .QN(n1244) );
  DFFRX1 \R_reg[11][2]  ( .D(n2277), .CK(clk), .RN(reset_n), .Q(\R[11][2] ), 
        .QN(n1243) );
  DFFRX1 \R_reg[11][3]  ( .D(n2276), .CK(clk), .RN(reset_n), .Q(\R[11][3] ), 
        .QN(n1242) );
  DFFRX1 \R_reg[11][4]  ( .D(n2275), .CK(clk), .RN(reset_n), .Q(\R[11][4] ), 
        .QN(n1241) );
  DFFRX1 \R_reg[11][5]  ( .D(n2274), .CK(clk), .RN(reset_n), .Q(\R[11][5] ), 
        .QN(n1240) );
  DFFRX1 \R_reg[11][6]  ( .D(n2273), .CK(clk), .RN(reset_n), .Q(\R[11][6] ), 
        .QN(n1239) );
  DFFRX1 \R_reg[15][0]  ( .D(n2151), .CK(clk), .RN(reset_n), .Q(\R[15][0] ), 
        .QN(n1117) );
  DFFRX1 \R_reg[15][1]  ( .D(n2150), .CK(clk), .RN(reset_n), .Q(\R[15][1] ), 
        .QN(n1116) );
  DFFRX1 \R_reg[15][2]  ( .D(n2149), .CK(clk), .RN(reset_n), .Q(\R[15][2] ), 
        .QN(n1115) );
  DFFRX1 \R_reg[15][3]  ( .D(n2148), .CK(clk), .RN(reset_n), .Q(\R[15][3] ), 
        .QN(n1114) );
  DFFRX1 \R_reg[15][4]  ( .D(n2147), .CK(clk), .RN(reset_n), .Q(\R[15][4] ), 
        .QN(n1113) );
  DFFRX1 \R_reg[15][5]  ( .D(n2146), .CK(clk), .RN(reset_n), .Q(\R[15][5] ), 
        .QN(n1112) );
  DFFRX1 \R_reg[15][6]  ( .D(n2145), .CK(clk), .RN(reset_n), .Q(\R[15][6] ), 
        .QN(n1111) );
  DFFRX1 \R_reg[19][0]  ( .D(n2023), .CK(clk), .RN(reset_n), .Q(\R[19][0] ), 
        .QN(n989) );
  DFFRX1 \R_reg[19][1]  ( .D(n2022), .CK(clk), .RN(reset_n), .Q(\R[19][1] ), 
        .QN(n988) );
  DFFRX1 \R_reg[19][2]  ( .D(n2021), .CK(clk), .RN(reset_n), .Q(\R[19][2] ), 
        .QN(n987) );
  DFFRX1 \R_reg[19][3]  ( .D(n2020), .CK(clk), .RN(reset_n), .Q(\R[19][3] ), 
        .QN(n986) );
  DFFRX1 \R_reg[19][4]  ( .D(n2019), .CK(clk), .RN(reset_n), .Q(\R[19][4] ), 
        .QN(n985) );
  DFFRX1 \R_reg[19][5]  ( .D(n2018), .CK(clk), .RN(reset_n), .Q(\R[19][5] ), 
        .QN(n984) );
  DFFRX1 \R_reg[19][6]  ( .D(n2017), .CK(clk), .RN(reset_n), .Q(\R[19][6] ), 
        .QN(n983) );
  DFFRX1 \R_reg[23][0]  ( .D(n1895), .CK(clk), .RN(reset_n), .Q(\R[23][0] ), 
        .QN(n861) );
  DFFRX1 \R_reg[23][1]  ( .D(n1894), .CK(clk), .RN(reset_n), .Q(\R[23][1] ), 
        .QN(n860) );
  DFFRX1 \R_reg[23][2]  ( .D(n1893), .CK(clk), .RN(reset_n), .Q(\R[23][2] ), 
        .QN(n859) );
  DFFRX1 \R_reg[23][3]  ( .D(n1892), .CK(clk), .RN(reset_n), .Q(\R[23][3] ), 
        .QN(n858) );
  DFFRX1 \R_reg[23][4]  ( .D(n1891), .CK(clk), .RN(reset_n), .Q(\R[23][4] ), 
        .QN(n857) );
  DFFRX1 \R_reg[23][5]  ( .D(n1890), .CK(clk), .RN(reset_n), .Q(\R[23][5] ), 
        .QN(n856) );
  DFFRX1 \R_reg[23][6]  ( .D(n1889), .CK(clk), .RN(reset_n), .Q(\R[23][6] ), 
        .QN(n855) );
  DFFRX1 \R_reg[27][0]  ( .D(n1767), .CK(clk), .RN(reset_n), .Q(\R[27][0] ), 
        .QN(n733) );
  DFFRX1 \R_reg[27][1]  ( .D(n1766), .CK(clk), .RN(reset_n), .Q(\R[27][1] ), 
        .QN(n732) );
  DFFRX1 \R_reg[27][2]  ( .D(n1765), .CK(clk), .RN(reset_n), .Q(\R[27][2] ), 
        .QN(n731) );
  DFFRX1 \R_reg[27][3]  ( .D(n1764), .CK(clk), .RN(reset_n), .Q(\R[27][3] ), 
        .QN(n730) );
  DFFRX1 \R_reg[27][4]  ( .D(n1763), .CK(clk), .RN(reset_n), .Q(\R[27][4] ), 
        .QN(n729) );
  DFFRX1 \R_reg[27][5]  ( .D(n1762), .CK(clk), .RN(reset_n), .Q(\R[27][5] ), 
        .QN(n728) );
  DFFRX1 \R_reg[27][6]  ( .D(n1761), .CK(clk), .RN(reset_n), .Q(\R[27][6] ), 
        .QN(n727) );
  DFFRX1 \R_reg[31][0]  ( .D(n1639), .CK(clk), .RN(reset_n), .Q(\R[31][0] ), 
        .QN(n605) );
  DFFRX1 \R_reg[31][1]  ( .D(n1638), .CK(clk), .RN(reset_n), .Q(\R[31][1] ), 
        .QN(n604) );
  DFFRX1 \R_reg[31][2]  ( .D(n1637), .CK(clk), .RN(reset_n), .Q(\R[31][2] ), 
        .QN(n603) );
  DFFRX1 \R_reg[31][3]  ( .D(n1636), .CK(clk), .RN(reset_n), .Q(\R[31][3] ), 
        .QN(n602) );
  DFFRX1 \R_reg[31][4]  ( .D(n1635), .CK(clk), .RN(reset_n), .Q(\R[31][4] ), 
        .QN(n601) );
  DFFRX1 \R_reg[31][5]  ( .D(n1634), .CK(clk), .RN(reset_n), .Q(\R[31][5] ), 
        .QN(n600) );
  DFFRX1 \R_reg[31][6]  ( .D(n1633), .CK(clk), .RN(reset_n), .Q(\R[31][6] ), 
        .QN(n599) );
  DFFRX1 \R_reg[5][0]  ( .D(n2471), .CK(clk), .RN(reset_n), .Q(\R[5][0] ), 
        .QN(n1437) );
  DFFRX1 \R_reg[5][2]  ( .D(n2469), .CK(clk), .RN(reset_n), .Q(\R[5][2] ), 
        .QN(n1435) );
  DFFRX1 \R_reg[5][3]  ( .D(n2468), .CK(clk), .RN(reset_n), .Q(\R[5][3] ), 
        .QN(n1434) );
  DFFRX1 \R_reg[5][4]  ( .D(n2467), .CK(clk), .RN(reset_n), .Q(\R[5][4] ), 
        .QN(n1433) );
  DFFRX1 \R_reg[5][5]  ( .D(n2466), .CK(clk), .RN(reset_n), .Q(\R[5][5] ), 
        .QN(n1432) );
  DFFRX1 \R_reg[5][6]  ( .D(n2465), .CK(clk), .RN(reset_n), .Q(\R[5][6] ), 
        .QN(n1431) );
  DFFRX1 \R_reg[9][0]  ( .D(n2343), .CK(clk), .RN(reset_n), .Q(\R[9][0] ), 
        .QN(n1309) );
  DFFRX1 \R_reg[9][2]  ( .D(n2341), .CK(clk), .RN(reset_n), .Q(\R[9][2] ), 
        .QN(n1307) );
  DFFRX1 \R_reg[9][3]  ( .D(n2340), .CK(clk), .RN(reset_n), .Q(\R[9][3] ), 
        .QN(n1306) );
  DFFRX1 \R_reg[9][4]  ( .D(n2339), .CK(clk), .RN(reset_n), .Q(\R[9][4] ), 
        .QN(n1305) );
  DFFRX1 \R_reg[9][5]  ( .D(n2338), .CK(clk), .RN(reset_n), .Q(\R[9][5] ), 
        .QN(n1304) );
  DFFRX1 \R_reg[9][6]  ( .D(n2337), .CK(clk), .RN(reset_n), .Q(\R[9][6] ), 
        .QN(n1303) );
  DFFRX1 \R_reg[13][0]  ( .D(n2215), .CK(clk), .RN(reset_n), .Q(\R[13][0] ), 
        .QN(n1181) );
  DFFRX1 \R_reg[13][1]  ( .D(n2214), .CK(clk), .RN(reset_n), .Q(\R[13][1] ), 
        .QN(n1180) );
  DFFRX1 \R_reg[13][2]  ( .D(n2213), .CK(clk), .RN(reset_n), .Q(\R[13][2] ), 
        .QN(n1179) );
  DFFRX1 \R_reg[13][3]  ( .D(n2212), .CK(clk), .RN(reset_n), .Q(\R[13][3] ), 
        .QN(n1178) );
  DFFRX1 \R_reg[13][4]  ( .D(n2211), .CK(clk), .RN(reset_n), .Q(\R[13][4] ), 
        .QN(n1177) );
  DFFRX1 \R_reg[13][5]  ( .D(n2210), .CK(clk), .RN(reset_n), .Q(\R[13][5] ), 
        .QN(n1176) );
  DFFRX1 \R_reg[13][6]  ( .D(n2209), .CK(clk), .RN(reset_n), .Q(\R[13][6] ), 
        .QN(n1175) );
  DFFRX1 \R_reg[17][0]  ( .D(n2087), .CK(clk), .RN(reset_n), .Q(\R[17][0] ), 
        .QN(n1053) );
  DFFRX1 \R_reg[17][2]  ( .D(n2085), .CK(clk), .RN(reset_n), .Q(\R[17][2] ), 
        .QN(n1051) );
  DFFRX1 \R_reg[17][3]  ( .D(n2084), .CK(clk), .RN(reset_n), .Q(\R[17][3] ), 
        .QN(n1050) );
  DFFRX1 \R_reg[17][4]  ( .D(n2083), .CK(clk), .RN(reset_n), .Q(\R[17][4] ), 
        .QN(n1049) );
  DFFRX1 \R_reg[17][5]  ( .D(n2082), .CK(clk), .RN(reset_n), .Q(\R[17][5] ), 
        .QN(n1048) );
  DFFRX1 \R_reg[17][6]  ( .D(n2081), .CK(clk), .RN(reset_n), .Q(\R[17][6] ), 
        .QN(n1047) );
  DFFRX1 \R_reg[21][0]  ( .D(n1959), .CK(clk), .RN(reset_n), .Q(\R[21][0] ), 
        .QN(n925) );
  DFFRX1 \R_reg[21][2]  ( .D(n1957), .CK(clk), .RN(reset_n), .Q(\R[21][2] ), 
        .QN(n923) );
  DFFRX1 \R_reg[21][3]  ( .D(n1956), .CK(clk), .RN(reset_n), .Q(\R[21][3] ), 
        .QN(n922) );
  DFFRX1 \R_reg[21][4]  ( .D(n1955), .CK(clk), .RN(reset_n), .Q(\R[21][4] ), 
        .QN(n921) );
  DFFRX1 \R_reg[21][5]  ( .D(n1954), .CK(clk), .RN(reset_n), .Q(\R[21][5] ), 
        .QN(n920) );
  DFFRX1 \R_reg[21][6]  ( .D(n1953), .CK(clk), .RN(reset_n), .Q(\R[21][6] ), 
        .QN(n919) );
  DFFRX1 \R_reg[25][0]  ( .D(n1831), .CK(clk), .RN(reset_n), .Q(\R[25][0] ), 
        .QN(n797) );
  DFFRX1 \R_reg[25][2]  ( .D(n1829), .CK(clk), .RN(reset_n), .Q(\R[25][2] ), 
        .QN(n795) );
  DFFRX1 \R_reg[25][3]  ( .D(n1828), .CK(clk), .RN(reset_n), .Q(\R[25][3] ), 
        .QN(n794) );
  DFFRX1 \R_reg[25][4]  ( .D(n1827), .CK(clk), .RN(reset_n), .Q(\R[25][4] ), 
        .QN(n793) );
  DFFRX1 \R_reg[25][5]  ( .D(n1826), .CK(clk), .RN(reset_n), .Q(\R[25][5] ), 
        .QN(n792) );
  DFFRX1 \R_reg[25][6]  ( .D(n1825), .CK(clk), .RN(reset_n), .Q(\R[25][6] ), 
        .QN(n791) );
  DFFRX1 \R_reg[29][0]  ( .D(n1703), .CK(clk), .RN(reset_n), .Q(\R[29][0] ), 
        .QN(n669) );
  DFFRX1 \R_reg[29][2]  ( .D(n1701), .CK(clk), .RN(reset_n), .Q(\R[29][2] ), 
        .QN(n667) );
  DFFRX1 \R_reg[29][3]  ( .D(n1700), .CK(clk), .RN(reset_n), .Q(\R[29][3] ), 
        .QN(n666) );
  DFFRX1 \R_reg[29][4]  ( .D(n1699), .CK(clk), .RN(reset_n), .Q(\R[29][4] ), 
        .QN(n665) );
  DFFRX1 \R_reg[29][5]  ( .D(n1698), .CK(clk), .RN(reset_n), .Q(\R[29][5] ), 
        .QN(n664) );
  DFFRX1 \R_reg[29][6]  ( .D(n1697), .CK(clk), .RN(reset_n), .Q(\R[29][6] ), 
        .QN(n663) );
  DFFRX1 \R_reg[4][0]  ( .D(n2503), .CK(clk), .RN(reset_n), .Q(\R[4][0] ), 
        .QN(n1469) );
  DFFRX1 \R_reg[4][1]  ( .D(n2502), .CK(clk), .RN(reset_n), .Q(\R[4][1] ), 
        .QN(n1468) );
  DFFRX1 \R_reg[4][2]  ( .D(n2501), .CK(clk), .RN(reset_n), .Q(\R[4][2] ), 
        .QN(n1467) );
  DFFRX1 \R_reg[4][3]  ( .D(n2500), .CK(clk), .RN(reset_n), .Q(\R[4][3] ), 
        .QN(n1466) );
  DFFRX1 \R_reg[4][4]  ( .D(n2499), .CK(clk), .RN(reset_n), .Q(\R[4][4] ), 
        .QN(n1465) );
  DFFRX1 \R_reg[4][5]  ( .D(n2498), .CK(clk), .RN(reset_n), .Q(\R[4][5] ), 
        .QN(n1464) );
  DFFRX1 \R_reg[4][6]  ( .D(n2497), .CK(clk), .RN(reset_n), .Q(\R[4][6] ), 
        .QN(n1463) );
  DFFRX1 \R_reg[8][0]  ( .D(n2375), .CK(clk), .RN(reset_n), .Q(\R[8][0] ), 
        .QN(n1341) );
  DFFRX1 \R_reg[8][2]  ( .D(n2373), .CK(clk), .RN(reset_n), .Q(\R[8][2] ), 
        .QN(n1339) );
  DFFRX1 \R_reg[8][3]  ( .D(n2372), .CK(clk), .RN(reset_n), .Q(\R[8][3] ), 
        .QN(n1338) );
  DFFRX1 \R_reg[8][4]  ( .D(n2371), .CK(clk), .RN(reset_n), .Q(\R[8][4] ), 
        .QN(n1337) );
  DFFRX1 \R_reg[8][5]  ( .D(n2370), .CK(clk), .RN(reset_n), .Q(\R[8][5] ), 
        .QN(n1336) );
  DFFRX1 \R_reg[8][6]  ( .D(n2369), .CK(clk), .RN(reset_n), .Q(\R[8][6] ), 
        .QN(n1335) );
  DFFRX1 \R_reg[12][0]  ( .D(n2247), .CK(clk), .RN(reset_n), .Q(\R[12][0] ), 
        .QN(n1213) );
  DFFRX1 \R_reg[12][1]  ( .D(n2246), .CK(clk), .RN(reset_n), .Q(\R[12][1] ), 
        .QN(n1212) );
  DFFRX1 \R_reg[12][2]  ( .D(n2245), .CK(clk), .RN(reset_n), .Q(\R[12][2] ), 
        .QN(n1211) );
  DFFRX1 \R_reg[12][3]  ( .D(n2244), .CK(clk), .RN(reset_n), .Q(\R[12][3] ), 
        .QN(n1210) );
  DFFRX1 \R_reg[12][4]  ( .D(n2243), .CK(clk), .RN(reset_n), .Q(\R[12][4] ), 
        .QN(n1209) );
  DFFRX1 \R_reg[12][5]  ( .D(n2242), .CK(clk), .RN(reset_n), .Q(\R[12][5] ), 
        .QN(n1208) );
  DFFRX1 \R_reg[12][6]  ( .D(n2241), .CK(clk), .RN(reset_n), .Q(\R[12][6] ), 
        .QN(n1207) );
  DFFRX1 \R_reg[16][0]  ( .D(n2119), .CK(clk), .RN(reset_n), .Q(\R[16][0] ), 
        .QN(n1085) );
  DFFRX1 \R_reg[16][2]  ( .D(n2117), .CK(clk), .RN(reset_n), .Q(\R[16][2] ), 
        .QN(n1083) );
  DFFRX1 \R_reg[16][3]  ( .D(n2116), .CK(clk), .RN(reset_n), .Q(\R[16][3] ), 
        .QN(n1082) );
  DFFRX1 \R_reg[16][4]  ( .D(n2115), .CK(clk), .RN(reset_n), .Q(\R[16][4] ), 
        .QN(n1081) );
  DFFRX1 \R_reg[16][5]  ( .D(n2114), .CK(clk), .RN(reset_n), .Q(\R[16][5] ), 
        .QN(n1080) );
  DFFRX1 \R_reg[16][6]  ( .D(n2113), .CK(clk), .RN(reset_n), .Q(\R[16][6] ), 
        .QN(n1079) );
  DFFRX1 \R_reg[20][0]  ( .D(n1991), .CK(clk), .RN(reset_n), .Q(\R[20][0] ), 
        .QN(n957) );
  DFFRX1 \R_reg[20][2]  ( .D(n1989), .CK(clk), .RN(reset_n), .Q(\R[20][2] ), 
        .QN(n955) );
  DFFRX1 \R_reg[20][3]  ( .D(n1988), .CK(clk), .RN(reset_n), .Q(\R[20][3] ), 
        .QN(n954) );
  DFFRX1 \R_reg[20][4]  ( .D(n1987), .CK(clk), .RN(reset_n), .Q(\R[20][4] ), 
        .QN(n953) );
  DFFRX1 \R_reg[20][5]  ( .D(n1986), .CK(clk), .RN(reset_n), .Q(\R[20][5] ), 
        .QN(n952) );
  DFFRX1 \R_reg[20][6]  ( .D(n1985), .CK(clk), .RN(reset_n), .Q(\R[20][6] ), 
        .QN(n951) );
  DFFRX1 \R_reg[24][0]  ( .D(n1863), .CK(clk), .RN(reset_n), .Q(\R[24][0] ), 
        .QN(n829) );
  DFFRX1 \R_reg[24][2]  ( .D(n1861), .CK(clk), .RN(reset_n), .Q(\R[24][2] ), 
        .QN(n827) );
  DFFRX1 \R_reg[24][3]  ( .D(n1860), .CK(clk), .RN(reset_n), .Q(\R[24][3] ), 
        .QN(n826) );
  DFFRX1 \R_reg[24][4]  ( .D(n1859), .CK(clk), .RN(reset_n), .Q(\R[24][4] ), 
        .QN(n825) );
  DFFRX1 \R_reg[24][5]  ( .D(n1858), .CK(clk), .RN(reset_n), .Q(\R[24][5] ), 
        .QN(n824) );
  DFFRX1 \R_reg[24][6]  ( .D(n1857), .CK(clk), .RN(reset_n), .Q(\R[24][6] ), 
        .QN(n823) );
  DFFRX1 \R_reg[28][0]  ( .D(n1735), .CK(clk), .RN(reset_n), .Q(\R[28][0] ), 
        .QN(n701) );
  DFFRX1 \R_reg[28][2]  ( .D(n1733), .CK(clk), .RN(reset_n), .Q(\R[28][2] ), 
        .QN(n699) );
  DFFRX1 \R_reg[28][3]  ( .D(n1732), .CK(clk), .RN(reset_n), .Q(\R[28][3] ), 
        .QN(n698) );
  DFFRX1 \R_reg[28][4]  ( .D(n1731), .CK(clk), .RN(reset_n), .Q(\R[28][4] ), 
        .QN(n697) );
  DFFRX1 \R_reg[28][5]  ( .D(n1730), .CK(clk), .RN(reset_n), .Q(\R[28][5] ), 
        .QN(n696) );
  DFFRX1 \R_reg[28][6]  ( .D(n1729), .CK(clk), .RN(reset_n), .Q(\R[28][6] ), 
        .QN(n695) );
  DFFRX1 \R_reg[6][0]  ( .D(n2439), .CK(clk), .RN(reset_n), .Q(\R[6][0] ), 
        .QN(n1405) );
  DFFRX1 \R_reg[6][1]  ( .D(n2438), .CK(clk), .RN(reset_n), .Q(\R[6][1] ), 
        .QN(n1404) );
  DFFRX1 \R_reg[6][2]  ( .D(n2437), .CK(clk), .RN(reset_n), .Q(\R[6][2] ), 
        .QN(n1403) );
  DFFRX1 \R_reg[6][3]  ( .D(n2436), .CK(clk), .RN(reset_n), .Q(\R[6][3] ), 
        .QN(n1402) );
  DFFRX1 \R_reg[6][4]  ( .D(n2435), .CK(clk), .RN(reset_n), .Q(\R[6][4] ), 
        .QN(n1401) );
  DFFRX1 \R_reg[6][5]  ( .D(n2434), .CK(clk), .RN(reset_n), .Q(\R[6][5] ), 
        .QN(n1400) );
  DFFRX1 \R_reg[6][6]  ( .D(n2433), .CK(clk), .RN(reset_n), .Q(\R[6][6] ), 
        .QN(n1399) );
  DFFRX1 \R_reg[10][0]  ( .D(n2311), .CK(clk), .RN(reset_n), .Q(\R[10][0] ), 
        .QN(n1277) );
  DFFRX1 \R_reg[10][1]  ( .D(n2310), .CK(clk), .RN(reset_n), .Q(\R[10][1] ), 
        .QN(n1276) );
  DFFRX1 \R_reg[10][2]  ( .D(n2309), .CK(clk), .RN(reset_n), .Q(\R[10][2] ), 
        .QN(n1275) );
  DFFRX1 \R_reg[10][3]  ( .D(n2308), .CK(clk), .RN(reset_n), .Q(\R[10][3] ), 
        .QN(n1274) );
  DFFRX1 \R_reg[10][4]  ( .D(n2307), .CK(clk), .RN(reset_n), .Q(\R[10][4] ), 
        .QN(n1273) );
  DFFRX1 \R_reg[10][5]  ( .D(n2306), .CK(clk), .RN(reset_n), .Q(\R[10][5] ), 
        .QN(n1272) );
  DFFRX1 \R_reg[10][6]  ( .D(n2305), .CK(clk), .RN(reset_n), .Q(\R[10][6] ), 
        .QN(n1271) );
  DFFRX1 \R_reg[14][0]  ( .D(n2183), .CK(clk), .RN(reset_n), .Q(\R[14][0] ), 
        .QN(n1149) );
  DFFRX1 \R_reg[14][1]  ( .D(n2182), .CK(clk), .RN(reset_n), .Q(\R[14][1] ), 
        .QN(n1148) );
  DFFRX1 \R_reg[14][2]  ( .D(n2181), .CK(clk), .RN(reset_n), .Q(\R[14][2] ), 
        .QN(n1147) );
  DFFRX1 \R_reg[14][3]  ( .D(n2180), .CK(clk), .RN(reset_n), .Q(\R[14][3] ), 
        .QN(n1146) );
  DFFRX1 \R_reg[14][4]  ( .D(n2179), .CK(clk), .RN(reset_n), .Q(\R[14][4] ), 
        .QN(n1145) );
  DFFRX1 \R_reg[14][5]  ( .D(n2178), .CK(clk), .RN(reset_n), .Q(\R[14][5] ), 
        .QN(n1144) );
  DFFRX1 \R_reg[14][6]  ( .D(n2177), .CK(clk), .RN(reset_n), .Q(\R[14][6] ), 
        .QN(n1143) );
  DFFRX1 \R_reg[18][0]  ( .D(n2055), .CK(clk), .RN(reset_n), .Q(\R[18][0] ), 
        .QN(n1021) );
  DFFRX1 \R_reg[18][1]  ( .D(n2054), .CK(clk), .RN(reset_n), .Q(\R[18][1] ), 
        .QN(n1020) );
  DFFRX1 \R_reg[18][2]  ( .D(n2053), .CK(clk), .RN(reset_n), .Q(\R[18][2] ), 
        .QN(n1019) );
  DFFRX1 \R_reg[18][3]  ( .D(n2052), .CK(clk), .RN(reset_n), .Q(\R[18][3] ), 
        .QN(n1018) );
  DFFRX1 \R_reg[18][4]  ( .D(n2051), .CK(clk), .RN(reset_n), .Q(\R[18][4] ), 
        .QN(n1017) );
  DFFRX1 \R_reg[18][5]  ( .D(n2050), .CK(clk), .RN(reset_n), .Q(\R[18][5] ), 
        .QN(n1016) );
  DFFRX1 \R_reg[18][6]  ( .D(n2049), .CK(clk), .RN(reset_n), .Q(\R[18][6] ), 
        .QN(n1015) );
  DFFRX1 \R_reg[22][0]  ( .D(n1927), .CK(clk), .RN(reset_n), .Q(\R[22][0] ), 
        .QN(n893) );
  DFFRX1 \R_reg[22][1]  ( .D(n1926), .CK(clk), .RN(reset_n), .Q(\R[22][1] ), 
        .QN(n892) );
  DFFRX1 \R_reg[22][2]  ( .D(n1925), .CK(clk), .RN(reset_n), .Q(\R[22][2] ), 
        .QN(n891) );
  DFFRX1 \R_reg[22][3]  ( .D(n1924), .CK(clk), .RN(reset_n), .Q(\R[22][3] ), 
        .QN(n890) );
  DFFRX1 \R_reg[22][4]  ( .D(n1923), .CK(clk), .RN(reset_n), .Q(\R[22][4] ), 
        .QN(n889) );
  DFFRX1 \R_reg[22][5]  ( .D(n1922), .CK(clk), .RN(reset_n), .Q(\R[22][5] ), 
        .QN(n888) );
  DFFRX1 \R_reg[22][6]  ( .D(n1921), .CK(clk), .RN(reset_n), .Q(\R[22][6] ), 
        .QN(n887) );
  DFFRX1 \R_reg[26][0]  ( .D(n1799), .CK(clk), .RN(reset_n), .Q(\R[26][0] ), 
        .QN(n765) );
  DFFRX1 \R_reg[26][1]  ( .D(n1798), .CK(clk), .RN(reset_n), .Q(\R[26][1] ), 
        .QN(n764) );
  DFFRX1 \R_reg[26][2]  ( .D(n1797), .CK(clk), .RN(reset_n), .Q(\R[26][2] ), 
        .QN(n763) );
  DFFRX1 \R_reg[26][3]  ( .D(n1796), .CK(clk), .RN(reset_n), .Q(\R[26][3] ), 
        .QN(n762) );
  DFFRX1 \R_reg[26][4]  ( .D(n1795), .CK(clk), .RN(reset_n), .Q(\R[26][4] ), 
        .QN(n761) );
  DFFRX1 \R_reg[26][5]  ( .D(n1794), .CK(clk), .RN(reset_n), .Q(\R[26][5] ), 
        .QN(n760) );
  DFFRX1 \R_reg[26][6]  ( .D(n1793), .CK(clk), .RN(reset_n), .Q(\R[26][6] ), 
        .QN(n759) );
  DFFRX1 \R_reg[30][0]  ( .D(n1671), .CK(clk), .RN(reset_n), .Q(\R[30][0] ), 
        .QN(n637) );
  DFFRX1 \R_reg[30][1]  ( .D(n1670), .CK(clk), .RN(reset_n), .Q(\R[30][1] ), 
        .QN(n636) );
  DFFRX1 \R_reg[30][2]  ( .D(n1669), .CK(clk), .RN(reset_n), .Q(\R[30][2] ), 
        .QN(n635) );
  DFFRX1 \R_reg[30][3]  ( .D(n1668), .CK(clk), .RN(reset_n), .Q(\R[30][3] ), 
        .QN(n634) );
  DFFRX1 \R_reg[30][4]  ( .D(n1667), .CK(clk), .RN(reset_n), .Q(\R[30][4] ), 
        .QN(n633) );
  DFFRX1 \R_reg[30][5]  ( .D(n1666), .CK(clk), .RN(reset_n), .Q(\R[30][5] ), 
        .QN(n632) );
  DFFRX1 \R_reg[30][6]  ( .D(n1665), .CK(clk), .RN(reset_n), .Q(\R[30][6] ), 
        .QN(n631) );
  DFFRX1 \R_reg[1][0]  ( .D(n2599), .CK(clk), .RN(reset_n), .Q(\R[1][0] ), 
        .QN(n1565) );
  DFFRX1 \R_reg[1][1]  ( .D(n2598), .CK(clk), .RN(reset_n), .Q(\R[1][1] ), 
        .QN(n1564) );
  DFFRX1 \R_reg[1][2]  ( .D(n2597), .CK(clk), .RN(reset_n), .Q(\R[1][2] ), 
        .QN(n1563) );
  DFFRX1 \R_reg[1][3]  ( .D(n2596), .CK(clk), .RN(reset_n), .Q(\R[1][3] ), 
        .QN(n1562) );
  DFFRX1 \R_reg[1][4]  ( .D(n2595), .CK(clk), .RN(reset_n), .Q(\R[1][4] ), 
        .QN(n1561) );
  DFFRX1 \R_reg[1][5]  ( .D(n2594), .CK(clk), .RN(reset_n), .Q(\R[1][5] ), 
        .QN(n1560) );
  DFFRX1 \R_reg[1][6]  ( .D(n2593), .CK(clk), .RN(reset_n), .Q(\R[1][6] ), 
        .QN(n1559) );
  DFFRX1 \R_reg[3][0]  ( .D(n2535), .CK(clk), .RN(reset_n), .Q(\R[3][0] ), 
        .QN(n1501) );
  DFFRX1 \R_reg[3][2]  ( .D(n2533), .CK(clk), .RN(reset_n), .Q(\R[3][2] ), 
        .QN(n1499) );
  DFFRX1 \R_reg[3][3]  ( .D(n2532), .CK(clk), .RN(reset_n), .Q(\R[3][3] ), 
        .QN(n1498) );
  DFFRX1 \R_reg[3][4]  ( .D(n2531), .CK(clk), .RN(reset_n), .Q(\R[3][4] ), 
        .QN(n1497) );
  DFFRX1 \R_reg[3][5]  ( .D(n2530), .CK(clk), .RN(reset_n), .Q(\R[3][5] ), 
        .QN(n1496) );
  DFFRX1 \R_reg[3][6]  ( .D(n2529), .CK(clk), .RN(reset_n), .Q(\R[3][6] ), 
        .QN(n1495) );
  DFFRX1 \R_reg[2][0]  ( .D(n2567), .CK(clk), .RN(reset_n), .QN(n1533) );
  DFFRX1 \R_reg[2][1]  ( .D(n2566), .CK(clk), .RN(reset_n), .QN(n1532) );
  DFFRX1 \R_reg[2][2]  ( .D(n2565), .CK(clk), .RN(reset_n), .QN(n1531) );
  DFFRX1 \R_reg[2][3]  ( .D(n2564), .CK(clk), .RN(reset_n), .QN(n1530) );
  DFFRX1 \R_reg[2][4]  ( .D(n2563), .CK(clk), .RN(reset_n), .QN(n1529) );
  DFFRX1 \R_reg[2][5]  ( .D(n2562), .CK(clk), .RN(reset_n), .QN(n1528) );
  DFFRX1 \R_reg[2][6]  ( .D(n2561), .CK(clk), .RN(reset_n), .QN(n1527) );
  DFFRX1 \R_reg[5][1]  ( .D(n2470), .CK(clk), .RN(reset_n), .Q(\R[5][1] ), 
        .QN(n1436) );
  DFFRX1 \R_reg[9][1]  ( .D(n2342), .CK(clk), .RN(reset_n), .Q(\R[9][1] ), 
        .QN(n1308) );
  DFFRX1 \R_reg[17][1]  ( .D(n2086), .CK(clk), .RN(reset_n), .Q(\R[17][1] ), 
        .QN(n1052) );
  DFFRX1 \R_reg[21][1]  ( .D(n1958), .CK(clk), .RN(reset_n), .Q(\R[21][1] ), 
        .QN(n924) );
  DFFRX1 \R_reg[25][1]  ( .D(n1830), .CK(clk), .RN(reset_n), .Q(\R[25][1] ), 
        .QN(n796) );
  DFFRX1 \R_reg[29][1]  ( .D(n1702), .CK(clk), .RN(reset_n), .Q(\R[29][1] ), 
        .QN(n668) );
  DFFRX1 \R_reg[8][1]  ( .D(n2374), .CK(clk), .RN(reset_n), .Q(\R[8][1] ), 
        .QN(n1340) );
  DFFRX1 \R_reg[16][1]  ( .D(n2118), .CK(clk), .RN(reset_n), .Q(\R[16][1] ), 
        .QN(n1084) );
  DFFRX1 \R_reg[20][1]  ( .D(n1990), .CK(clk), .RN(reset_n), .Q(\R[20][1] ), 
        .QN(n956) );
  DFFRX1 \R_reg[24][1]  ( .D(n1862), .CK(clk), .RN(reset_n), .Q(\R[24][1] ), 
        .QN(n828) );
  DFFRX1 \R_reg[28][1]  ( .D(n1734), .CK(clk), .RN(reset_n), .Q(\R[28][1] ), 
        .QN(n700) );
  DFFRX1 \R_reg[3][1]  ( .D(n2534), .CK(clk), .RN(reset_n), .Q(\R[3][1] ), 
        .QN(n1500) );
  DFFRX1 \R_reg[10][31]  ( .D(n2280), .CK(clk), .RN(reset_n), .Q(\R[10][31] )
         );
  MXI2X2 U1694 ( .A(n2681), .B(n2682), .S0(n3231), .Y(n2663) );
  MX4X2 U1695 ( .A(n2761), .B(n2762), .C(n2763), .D(n2764), .S0(n3223), .S1(
        n3215), .Y(n2682) );
  MXI2X4 U1696 ( .A(n2681), .B(n2682), .S0(n3231), .Y(n2670) );
  XOR2X1 U1697 ( .A(n4043), .B(\sub_1_root_add_0_root_add_137_ni_b0/carry[6] ), 
        .Y(N650) );
  NAND2X1 U1698 ( .A(n2662), .B(n3215), .Y(n2660) );
  CLKMX2X2 U1699 ( .A(n3270), .B(n3265), .S0(n3767), .Y(N250) );
  MXI4X1 U1700 ( .A(n3291), .B(n3292), .C(n3293), .D(n3294), .S0(n3760), .S1(
        n3752), .Y(n3290) );
  MX4X1 U1701 ( .A(n2769), .B(n2770), .C(n2771), .D(n2772), .S0(n3223), .S1(
        n3215), .Y(n2680) );
  MXI2X2 U1702 ( .A(n2748), .B(n2749), .S0(n3232), .Y(n2673) );
  MXI4X1 U1703 ( .A(\R[24][10] ), .B(\R[25][10] ), .C(\R[26][10] ), .D(
        \R[27][10] ), .S0(n3180), .S1(n3207), .Y(n2842) );
  MXI2X2 U1704 ( .A(n2753), .B(n2754), .S0(n3232), .Y(n2674) );
  MXI2X1 U1705 ( .A(n2755), .B(n2756), .S0(n3232), .Y(n2675) );
  MX4X1 U1706 ( .A(n2825), .B(n2826), .C(n2827), .D(n2828), .S0(n3225), .S1(
        n3217), .Y(n2756) );
  MXI2X2 U1707 ( .A(n2757), .B(n2758), .S0(n3231), .Y(n2671) );
  MX4X1 U1708 ( .A(n2817), .B(n2818), .C(n2819), .D(n2820), .S0(n3224), .S1(
        n3216), .Y(n2758) );
  MXI2X2 U1709 ( .A(n2691), .B(n2692), .S0(n3231), .Y(n2672) );
  MX4X1 U1710 ( .A(n2805), .B(n2806), .C(n2807), .D(n2808), .S0(n3224), .S1(
        n3216), .Y(n2689) );
  MXI4X1 U1711 ( .A(\R[24][5] ), .B(\R[25][5] ), .C(\R[26][5] ), .D(\R[27][5] ), .S0(n3179), .S1(n3207), .Y(n2802) );
  MXI2X2 U1712 ( .A(n2744), .B(n2745), .S0(n3232), .Y(n2677) );
  AND4X1 U1713 ( .A(n325), .B(n326), .C(n327), .D(n328), .Y(n125) );
  AND4X1 U1714 ( .A(n331), .B(n332), .C(n333), .D(n334), .Y(n126) );
  MX4X1 U1715 ( .A(n2793), .B(n2794), .C(n2795), .D(n2796), .S0(n3224), .S1(
        n3216), .Y(n2688) );
  MX4X1 U1716 ( .A(n2797), .B(n2798), .C(n2799), .D(n2800), .S0(n3224), .S1(
        n3216), .Y(n2687) );
  MXI4X1 U1717 ( .A(\R[24][4] ), .B(\R[25][4] ), .C(\R[26][4] ), .D(\R[27][4] ), .S0(n3179), .S1(n3207), .Y(n2794) );
  CLKBUFX3 U1718 ( .A(n130), .Y(n3919) );
  MXI2X2 U1719 ( .A(n2702), .B(n2703), .S0(n3233), .Y(n2648) );
  MXI2X2 U1720 ( .A(n2731), .B(n2732), .S0(n3232), .Y(n2649) );
  MXI2X2 U1721 ( .A(n2723), .B(n2724), .S0(n3233), .Y(n2650) );
  MXI2X2 U1722 ( .A(n2721), .B(n2722), .S0(n3233), .Y(n2651) );
  MXI2X2 U1723 ( .A(n2719), .B(n2720), .S0(n3233), .Y(n2652) );
  MXI2X2 U1724 ( .A(n2733), .B(n2734), .S0(n3232), .Y(n2653) );
  CLKINVX1 U1725 ( .A(n2707), .Y(N199) );
  INVX1 U1726 ( .A(n2693), .Y(N218) );
  CLKMX2X2 U1727 ( .A(n2694), .B(n2695), .S0(n3231), .Y(n2693) );
  NOR2X1 U1728 ( .A(n3992), .B(n3991), .Y(n2654) );
  MXI2X2 U1729 ( .A(n2689), .B(n2690), .S0(n3231), .Y(n2655) );
  CLKINVX1 U1730 ( .A(n2725), .Y(N198) );
  INVX1 U1731 ( .A(n2683), .Y(N219) );
  CLKMX2X2 U1732 ( .A(n2684), .B(n2685), .S0(n3231), .Y(n2683) );
  CLKINVX1 U1733 ( .A(n2686), .Y(N217) );
  CLKMX2X2 U1734 ( .A(n2687), .B(n2688), .S0(n3231), .Y(n2686) );
  NOR2X1 U1735 ( .A(n3998), .B(n243), .Y(n2656) );
  NOR2X2 U1736 ( .A(\sub_1_root_add_0_root_add_137_ni_b0/carry[14] ), .B(
        \seIM[31] ), .Y(n2657) );
  AND4X4 U1737 ( .A(n311), .B(n312), .C(n313), .D(n314), .Y(n123) );
  AOI222X1 U1738 ( .A0(N926), .A1(n3777), .B0(N894), .B1(n251), .C0(N815), 
        .C1(n249), .Y(n312) );
  MX4X1 U1739 ( .A(n2841), .B(n2842), .C(n2843), .D(n2844), .S0(n3225), .S1(
        n3217), .Y(n2749) );
  CLKBUFX3 U1740 ( .A(n3221), .Y(n3215) );
  NAND2X1 U1741 ( .A(n2661), .B(n2658), .Y(n2659) );
  NAND2X2 U1742 ( .A(n2659), .B(n2660), .Y(n2681) );
  INVXL U1743 ( .A(n3215), .Y(n2658) );
  CLKINVX1 U1744 ( .A(n2750), .Y(N207) );
  MXI4XL U1745 ( .A(\R[12][3] ), .B(\R[13][3] ), .C(\R[14][3] ), .D(\R[15][3] ), .S0(n3717), .S1(n3742), .Y(n3274) );
  CLKMX2X2 U1746 ( .A(n3380), .B(n3375), .S0(n3768), .Y(N239) );
  INVX4 U1747 ( .A(n2678), .Y(N220) );
  CLKBUFX3 U1748 ( .A(n3229), .Y(n3223) );
  MX2X2 U1749 ( .A(n2765), .B(n2766), .S0(n3223), .Y(n2661) );
  MX2X2 U1750 ( .A(n2767), .B(n2768), .S0(n3223), .Y(n2662) );
  CLKBUFX2 U1751 ( .A(n131), .Y(n3915) );
  CLKBUFX2 U1752 ( .A(n131), .Y(n3914) );
  AOI222X1 U1753 ( .A0(N688), .A1(n247), .B0(N190), .B1(n307), .C0(N222), .C1(
        n308), .Y(n306) );
  NOR2X1 U1754 ( .A(n2669), .B(n2667), .Y(n2664) );
  NOR2X1 U1755 ( .A(n2665), .B(n2668), .Y(n305) );
  CLKINVX1 U1756 ( .A(n2664), .Y(n2665) );
  AND2X2 U1757 ( .A(N464), .B(n246), .Y(n2669) );
  CLKBUFX2 U1758 ( .A(n122), .Y(n3943) );
  MX2X2 U1759 ( .A(n2679), .B(n2680), .S0(n3231), .Y(n2678) );
  BUFX2 U1760 ( .A(n131), .Y(n3916) );
  AOI222XL U1761 ( .A0(N924), .A1(n3777), .B0(N892), .B1(n251), .C0(N813), 
        .C1(n249), .Y(n332) );
  OAI2BB2XL U1762 ( .B0(n3943), .B1(n3796), .A0N(\R[10][31] ), .A1N(n3794), 
        .Y(n2280) );
  CLKBUFX3 U1763 ( .A(n130), .Y(n3918) );
  CLKBUFX3 U1764 ( .A(n130), .Y(n3917) );
  CLKBUFX3 U1765 ( .A(n132), .Y(n3911) );
  CLKBUFX3 U1766 ( .A(n132), .Y(n3913) );
  AND2X2 U1767 ( .A(n551), .B(n524), .Y(n3780) );
  OAI22XL U1768 ( .A0(n1248), .A1(n3798), .B0(n3934), .B1(n3796), .Y(n2282) );
  AOI222X1 U1769 ( .A0(N927), .A1(n253), .B0(N895), .B1(n3778), .C0(N816), 
        .C1(n249), .Y(n304) );
  OAI22XL U1770 ( .A0(n1249), .A1(n3798), .B0(n3931), .B1(n3796), .Y(n2283) );
  OAI22XL U1771 ( .A0(n1250), .A1(n3798), .B0(n3928), .B1(n3796), .Y(n2284) );
  OAI22XL U1772 ( .A0(n1251), .A1(n3798), .B0(n3925), .B1(n3796), .Y(n2285) );
  OAI22XL U1773 ( .A0(n1252), .A1(n3798), .B0(n3922), .B1(n3796), .Y(n2286) );
  MXI4XL U1774 ( .A(\R[12][5] ), .B(\R[13][5] ), .C(\R[14][5] ), .D(\R[15][5] ), .S0(n3717), .S1(n3743), .Y(n3294) );
  CLKMX2X2 U1775 ( .A(n3290), .B(n3285), .S0(n3767), .Y(N248) );
  MXI4X1 U1776 ( .A(\R[20][12] ), .B(\R[21][12] ), .C(\R[22][12] ), .D(
        \R[23][12] ), .S0(n3180), .S1(n3207), .Y(n2859) );
  MXI4X1 U1777 ( .A(\R[4][12] ), .B(\R[5][12] ), .C(\R[6][12] ), .D(\R[7][12] ), .S0(n3180), .S1(n3207), .Y(n2863) );
  MXI4X1 U1778 ( .A(\R[24][12] ), .B(\R[25][12] ), .C(\R[26][12] ), .D(
        \R[27][12] ), .S0(n3180), .S1(n3207), .Y(n2858) );
  MXI4X1 U1779 ( .A(\R[8][12] ), .B(\R[9][12] ), .C(\R[10][12] ), .D(
        \R[11][12] ), .S0(n3180), .S1(n3207), .Y(n2862) );
  MXI4X1 U1780 ( .A(\R[24][11] ), .B(\R[25][11] ), .C(\R[26][11] ), .D(
        \R[27][11] ), .S0(n3180), .S1(n3207), .Y(n2850) );
  MXI4X1 U1781 ( .A(\R[8][11] ), .B(\R[9][11] ), .C(\R[10][11] ), .D(
        \R[11][11] ), .S0(n3180), .S1(n3207), .Y(n2854) );
  INVXL U1782 ( .A(N220), .Y(n4023) );
  AND2X2 U1783 ( .A(N432), .B(n3779), .Y(n2667) );
  AND2X2 U1784 ( .A(N624), .B(n3780), .Y(n2668) );
  AND2XL U1785 ( .A(n562), .B(n553), .Y(n246) );
  AND4X4 U1786 ( .A(n306), .B(n304), .C(n305), .D(n303), .Y(n122) );
  CLKBUFX3 U1787 ( .A(n3187), .Y(n3181) );
  MX4X2 U1788 ( .A(n2781), .B(n2782), .C(n2783), .D(n2784), .S0(n3224), .S1(
        n3216), .Y(n2684) );
  MX4X2 U1789 ( .A(n2777), .B(n2778), .C(n2779), .D(n2780), .S0(n3224), .S1(
        n3216), .Y(n2685) );
  MX4X2 U1790 ( .A(n2789), .B(n2790), .C(n2791), .D(n2792), .S0(n3224), .S1(
        n3216), .Y(n2694) );
  MX4X2 U1791 ( .A(n2785), .B(n2786), .C(n2787), .D(n2788), .S0(n3224), .S1(
        n3216), .Y(n2695) );
  CLKBUFX2 U1792 ( .A(n127), .Y(n3928) );
  CLKBUFX2 U1793 ( .A(n128), .Y(n3925) );
  CLKBUFX2 U1794 ( .A(n129), .Y(n3922) );
  BUFX2 U1795 ( .A(n132), .Y(n3912) );
  MXI2X2 U1796 ( .A(n2746), .B(n2747), .S0(n3232), .Y(n2676) );
  CLKINVX1 U1797 ( .A(n465), .Y(n4045) );
  INVXL U1798 ( .A(N241), .Y(n4027) );
  INVXL U1799 ( .A(N243), .Y(n4029) );
  INVXL U1800 ( .A(N245), .Y(n4031) );
  INVXL U1801 ( .A(N246), .Y(n4032) );
  INVXL U1802 ( .A(N249), .Y(n4035) );
  INVXL U1803 ( .A(N242), .Y(n4028) );
  INVXL U1804 ( .A(N244), .Y(n4030) );
  INVXL U1805 ( .A(N252), .Y(n4038) );
  INVXL U1806 ( .A(N247), .Y(n4033) );
  INVXL U1807 ( .A(N250), .Y(n4036) );
  INVXL U1808 ( .A(N251), .Y(n4037) );
  INVXL U1809 ( .A(N253), .Y(n4039) );
  NAND2X1 U1810 ( .A(n561), .B(n560), .Y(n237) );
  CLKINVX1 U1811 ( .A(n3981), .Y(n3980) );
  OAI22X1 U1812 ( .A0(n1247), .A1(n3798), .B0(n3940), .B1(n3796), .Y(n2281) );
  NOR2XL U1813 ( .A(n3750), .B(\R[1][1] ), .Y(n3707) );
  NOR2XL U1814 ( .A(n3750), .B(\R[1][0] ), .Y(n3712) );
  NOR2XL U1815 ( .A(\R[3][1] ), .B(n3740), .Y(n3705) );
  NOR2XL U1816 ( .A(\R[3][0] ), .B(n3741), .Y(n3710) );
  MXI4XL U1817 ( .A(\R[28][1] ), .B(\R[29][1] ), .C(\R[30][1] ), .D(\R[31][1] ), .S0(n3717), .S1(n3742), .Y(n3249) );
  MXI4XL U1818 ( .A(\R[12][0] ), .B(\R[13][0] ), .C(\R[14][0] ), .D(\R[15][0] ), .S0(n3717), .S1(n3742), .Y(n3244) );
  MXI4XL U1819 ( .A(\R[20][1] ), .B(\R[21][1] ), .C(\R[22][1] ), .D(\R[23][1] ), .S0(n3717), .S1(n3742), .Y(n3248) );
  MXI4XL U1820 ( .A(\R[4][1] ), .B(\R[5][1] ), .C(\R[6][1] ), .D(\R[7][1] ), 
        .S0(n3717), .S1(n3742), .Y(n3253) );
  MXI4XL U1821 ( .A(\R[4][0] ), .B(\R[5][0] ), .C(\R[6][0] ), .D(\R[7][0] ), 
        .S0(n3717), .S1(n3742), .Y(n3243) );
  MXI4XL U1822 ( .A(\R[20][0] ), .B(\R[21][0] ), .C(\R[22][0] ), .D(\R[23][0] ), .S0(n3717), .S1(n3742), .Y(n3238) );
  MXI4XL U1823 ( .A(\R[16][1] ), .B(\R[17][1] ), .C(\R[18][1] ), .D(\R[19][1] ), .S0(n3717), .S1(n3742), .Y(n3246) );
  MXI4XL U1824 ( .A(\R[16][0] ), .B(\R[17][0] ), .C(\R[18][0] ), .D(\R[19][0] ), .S0(n3717), .S1(n3742), .Y(n3236) );
  MXI4XL U1825 ( .A(\R[8][1] ), .B(\R[9][1] ), .C(\R[10][1] ), .D(\R[11][1] ), 
        .S0(n3717), .S1(n3742), .Y(n3252) );
  MXI4XL U1826 ( .A(\R[24][1] ), .B(\R[25][1] ), .C(\R[26][1] ), .D(\R[27][1] ), .S0(n3717), .S1(n3742), .Y(n3247) );
  MXI4XL U1827 ( .A(\R[8][0] ), .B(\R[9][0] ), .C(\R[10][0] ), .D(\R[11][0] ), 
        .S0(n3717), .S1(n3742), .Y(n3242) );
  MXI4XL U1828 ( .A(\R[24][0] ), .B(\R[25][0] ), .C(\R[26][0] ), .D(\R[27][0] ), .S0(n3717), .S1(n3742), .Y(n3237) );
  NOR2XL U1829 ( .A(n3750), .B(\R[1][2] ), .Y(n3702) );
  NOR2XL U1830 ( .A(n3750), .B(\R[1][3] ), .Y(n3697) );
  NOR2XL U1831 ( .A(n3750), .B(\R[1][4] ), .Y(n3692) );
  NOR2XL U1832 ( .A(\R[3][2] ), .B(n3739), .Y(n3700) );
  NOR2XL U1833 ( .A(\R[3][3] ), .B(n3738), .Y(n3695) );
  NOR2XL U1834 ( .A(\R[3][4] ), .B(n3737), .Y(n3690) );
  MXI4X2 U1835 ( .A(\R[8][4] ), .B(\R[9][4] ), .C(\R[10][4] ), .D(\R[11][4] ), 
        .S0(n3179), .S1(n3207), .Y(n2798) );
  MXI4XL U1836 ( .A(\R[28][2] ), .B(\R[29][2] ), .C(\R[30][2] ), .D(\R[31][2] ), .S0(n3717), .S1(n3742), .Y(n3259) );
  MXI4XL U1837 ( .A(\R[28][3] ), .B(\R[29][3] ), .C(\R[30][3] ), .D(\R[31][3] ), .S0(n3717), .S1(n3742), .Y(n3269) );
  MXI4XL U1838 ( .A(\R[28][4] ), .B(\R[29][4] ), .C(\R[30][4] ), .D(\R[31][4] ), .S0(n3717), .S1(n3743), .Y(n3279) );
  MXI4XL U1839 ( .A(\R[20][2] ), .B(\R[21][2] ), .C(\R[22][2] ), .D(\R[23][2] ), .S0(n3717), .S1(n3742), .Y(n3258) );
  MXI4XL U1840 ( .A(\R[4][2] ), .B(\R[5][2] ), .C(\R[6][2] ), .D(\R[7][2] ), 
        .S0(n3717), .S1(n3742), .Y(n3263) );
  MXI4XL U1841 ( .A(\R[20][3] ), .B(\R[21][3] ), .C(\R[22][3] ), .D(\R[23][3] ), .S0(n3717), .S1(n3742), .Y(n3268) );
  MXI4XL U1842 ( .A(\R[4][3] ), .B(\R[5][3] ), .C(\R[6][3] ), .D(\R[7][3] ), 
        .S0(n3717), .S1(n3742), .Y(n3273) );
  MXI4XL U1843 ( .A(\R[20][4] ), .B(\R[21][4] ), .C(\R[22][4] ), .D(\R[23][4] ), .S0(n3717), .S1(n3743), .Y(n3278) );
  MXI4XL U1844 ( .A(\R[4][4] ), .B(\R[5][4] ), .C(\R[6][4] ), .D(\R[7][4] ), 
        .S0(n3717), .S1(n3743), .Y(n3283) );
  MXI4XL U1845 ( .A(\R[16][2] ), .B(\R[17][2] ), .C(\R[18][2] ), .D(\R[19][2] ), .S0(n3717), .S1(n3742), .Y(n3256) );
  MXI4XL U1846 ( .A(\R[16][3] ), .B(\R[17][3] ), .C(\R[18][3] ), .D(\R[19][3] ), .S0(n3717), .S1(n3742), .Y(n3266) );
  MXI4XL U1847 ( .A(\R[16][4] ), .B(\R[17][4] ), .C(\R[18][4] ), .D(\R[19][4] ), .S0(n3717), .S1(n3743), .Y(n3276) );
  MXI4XL U1848 ( .A(\R[8][2] ), .B(\R[9][2] ), .C(\R[10][2] ), .D(\R[11][2] ), 
        .S0(n3717), .S1(n3742), .Y(n3262) );
  MXI4XL U1849 ( .A(\R[24][2] ), .B(\R[25][2] ), .C(\R[26][2] ), .D(\R[27][2] ), .S0(n3717), .S1(n3742), .Y(n3257) );
  MXI4XL U1850 ( .A(\R[8][3] ), .B(\R[9][3] ), .C(\R[10][3] ), .D(\R[11][3] ), 
        .S0(n3717), .S1(n3742), .Y(n3272) );
  MXI4XL U1851 ( .A(\R[24][3] ), .B(\R[25][3] ), .C(\R[26][3] ), .D(\R[27][3] ), .S0(n3717), .S1(n3742), .Y(n3267) );
  MXI4XL U1852 ( .A(\R[8][4] ), .B(\R[9][4] ), .C(\R[10][4] ), .D(\R[11][4] ), 
        .S0(n3717), .S1(n3743), .Y(n3282) );
  MXI4XL U1853 ( .A(\R[24][4] ), .B(\R[25][4] ), .C(\R[26][4] ), .D(\R[27][4] ), .S0(n3717), .S1(n3743), .Y(n3277) );
  AOI22XL U1854 ( .A0(N284), .A1(n3789), .B0(N1023), .B1(n3785), .Y(n489) );
  NOR2XL U1855 ( .A(n3750), .B(\R[1][5] ), .Y(n3687) );
  NOR2XL U1856 ( .A(n3750), .B(\R[1][6] ), .Y(n3682) );
  NOR2XL U1857 ( .A(\R[3][5] ), .B(n3736), .Y(n3685) );
  NOR2XL U1858 ( .A(\R[3][6] ), .B(n3735), .Y(n3680) );
  MXI4X2 U1859 ( .A(\R[12][5] ), .B(\R[13][5] ), .C(\R[14][5] ), .D(\R[15][5] ), .S0(n3179), .S1(n3207), .Y(n2808) );
  MXI4X2 U1860 ( .A(\R[28][5] ), .B(\R[29][5] ), .C(\R[30][5] ), .D(\R[31][5] ), .S0(n3179), .S1(n3207), .Y(n2804) );
  MXI4X2 U1861 ( .A(\R[16][5] ), .B(\R[17][5] ), .C(\R[18][5] ), .D(\R[19][5] ), .S0(n3179), .S1(n3207), .Y(n2801) );
  MXI4X2 U1862 ( .A(\R[20][5] ), .B(\R[21][5] ), .C(\R[22][5] ), .D(\R[23][5] ), .S0(n3179), .S1(n3207), .Y(n2803) );
  MXI4XL U1863 ( .A(\R[28][5] ), .B(\R[29][5] ), .C(\R[30][5] ), .D(\R[31][5] ), .S0(n3717), .S1(n3743), .Y(n3289) );
  MXI4XL U1864 ( .A(\R[28][6] ), .B(\R[29][6] ), .C(\R[30][6] ), .D(\R[31][6] ), .S0(n3718), .S1(n3743), .Y(n3299) );
  MXI4XL U1865 ( .A(\R[20][5] ), .B(\R[21][5] ), .C(\R[22][5] ), .D(\R[23][5] ), .S0(n3717), .S1(n3743), .Y(n3288) );
  MXI4XL U1866 ( .A(\R[4][5] ), .B(\R[5][5] ), .C(\R[6][5] ), .D(\R[7][5] ), 
        .S0(n3718), .S1(n3743), .Y(n3293) );
  MXI4XL U1867 ( .A(\R[20][6] ), .B(\R[21][6] ), .C(\R[22][6] ), .D(\R[23][6] ), .S0(n3718), .S1(n3743), .Y(n3298) );
  MXI4XL U1868 ( .A(\R[4][6] ), .B(\R[5][6] ), .C(\R[6][6] ), .D(\R[7][6] ), 
        .S0(n3718), .S1(n3743), .Y(n3303) );
  MXI4XL U1869 ( .A(\R[16][5] ), .B(\R[17][5] ), .C(\R[18][5] ), .D(\R[19][5] ), .S0(n3717), .S1(n3743), .Y(n3286) );
  MXI4XL U1870 ( .A(\R[16][6] ), .B(\R[17][6] ), .C(\R[18][6] ), .D(\R[19][6] ), .S0(n3718), .S1(n3743), .Y(n3296) );
  MXI4XL U1871 ( .A(\R[8][5] ), .B(\R[9][5] ), .C(\R[10][5] ), .D(\R[11][5] ), 
        .S0(n3718), .S1(n3743), .Y(n3292) );
  MXI4XL U1872 ( .A(\R[24][5] ), .B(\R[25][5] ), .C(\R[26][5] ), .D(\R[27][5] ), .S0(n3717), .S1(n3743), .Y(n3287) );
  MXI4XL U1873 ( .A(\R[8][6] ), .B(\R[9][6] ), .C(\R[10][6] ), .D(\R[11][6] ), 
        .S0(n3718), .S1(n3743), .Y(n3302) );
  MXI4XL U1874 ( .A(\R[24][6] ), .B(\R[25][6] ), .C(\R[26][6] ), .D(\R[27][6] ), .S0(n3718), .S1(n3743), .Y(n3297) );
  AOI22XL U1875 ( .A0(N282), .A1(n3789), .B0(N1021), .B1(n3785), .Y(n492) );
  AOI22XL U1876 ( .A0(N281), .A1(n3789), .B0(N1020), .B1(n3785), .Y(n493) );
  NOR2XL U1877 ( .A(n3749), .B(\R[1][7] ), .Y(n3677) );
  NOR2XL U1878 ( .A(n3749), .B(\R[1][8] ), .Y(n3672) );
  NOR2XL U1879 ( .A(n3749), .B(\R[1][9] ), .Y(n3667) );
  NOR2XL U1880 ( .A(\R[3][9] ), .B(n3732), .Y(n3665) );
  NOR2XL U1881 ( .A(\R[3][7] ), .B(n3734), .Y(n3675) );
  NOR2XL U1882 ( .A(\R[3][8] ), .B(n3733), .Y(n3670) );
  MXI4XL U1883 ( .A(\R[28][9] ), .B(\R[29][9] ), .C(\R[30][9] ), .D(\R[31][9] ), .S0(n3718), .S1(n3743), .Y(n3329) );
  MXI4XL U1884 ( .A(\R[28][8] ), .B(\R[29][8] ), .C(\R[30][8] ), .D(\R[31][8] ), .S0(n3718), .S1(n3743), .Y(n3319) );
  MXI4XL U1885 ( .A(\R[28][7] ), .B(\R[29][7] ), .C(\R[30][7] ), .D(\R[31][7] ), .S0(n3718), .S1(n3743), .Y(n3309) );
  MXI4XL U1886 ( .A(\R[20][9] ), .B(\R[21][9] ), .C(\R[22][9] ), .D(\R[23][9] ), .S0(n3718), .S1(n3743), .Y(n3328) );
  MXI4XL U1887 ( .A(\R[4][9] ), .B(\R[5][9] ), .C(\R[6][9] ), .D(\R[7][9] ), 
        .S0(n3718), .S1(n3743), .Y(n3333) );
  MXI4XL U1888 ( .A(\R[20][8] ), .B(\R[21][8] ), .C(\R[22][8] ), .D(\R[23][8] ), .S0(n3718), .S1(n3743), .Y(n3318) );
  MXI4XL U1889 ( .A(\R[4][8] ), .B(\R[5][8] ), .C(\R[6][8] ), .D(\R[7][8] ), 
        .S0(n3718), .S1(n3743), .Y(n3323) );
  MXI4XL U1890 ( .A(\R[20][7] ), .B(\R[21][7] ), .C(\R[22][7] ), .D(\R[23][7] ), .S0(n3718), .S1(n3743), .Y(n3308) );
  MXI4XL U1891 ( .A(\R[4][7] ), .B(\R[5][7] ), .C(\R[6][7] ), .D(\R[7][7] ), 
        .S0(n3718), .S1(n3743), .Y(n3313) );
  MXI4XL U1892 ( .A(\R[16][9] ), .B(\R[17][9] ), .C(\R[18][9] ), .D(\R[19][9] ), .S0(n3718), .S1(n3743), .Y(n3326) );
  MXI4XL U1893 ( .A(\R[16][8] ), .B(\R[17][8] ), .C(\R[18][8] ), .D(\R[19][8] ), .S0(n3718), .S1(n3743), .Y(n3316) );
  MXI4XL U1894 ( .A(\R[16][7] ), .B(\R[17][7] ), .C(\R[18][7] ), .D(\R[19][7] ), .S0(n3718), .S1(n3743), .Y(n3306) );
  MXI4XL U1895 ( .A(\R[8][9] ), .B(\R[9][9] ), .C(\R[10][9] ), .D(\R[11][9] ), 
        .S0(n3718), .S1(n3743), .Y(n3332) );
  MXI4XL U1896 ( .A(\R[24][9] ), .B(\R[25][9] ), .C(\R[26][9] ), .D(\R[27][9] ), .S0(n3718), .S1(n3743), .Y(n3327) );
  MXI4XL U1897 ( .A(\R[8][8] ), .B(\R[9][8] ), .C(\R[10][8] ), .D(\R[11][8] ), 
        .S0(n3718), .S1(n3743), .Y(n3322) );
  MXI4XL U1898 ( .A(\R[8][7] ), .B(\R[9][7] ), .C(\R[10][7] ), .D(\R[11][7] ), 
        .S0(n3718), .S1(n3743), .Y(n3312) );
  MXI4XL U1899 ( .A(\R[24][8] ), .B(\R[25][8] ), .C(\R[26][8] ), .D(\R[27][8] ), .S0(n3718), .S1(n3743), .Y(n3317) );
  MXI4XL U1900 ( .A(\R[24][7] ), .B(\R[25][7] ), .C(\R[26][7] ), .D(\R[27][7] ), .S0(n3718), .S1(n3743), .Y(n3307) );
  AOI22XL U1901 ( .A0(N280), .A1(n3789), .B0(N1019), .B1(n3785), .Y(n494) );
  AOI22XL U1902 ( .A0(N279), .A1(n3789), .B0(N1018), .B1(n3785), .Y(n495) );
  AOI22XL U1903 ( .A0(N278), .A1(n3789), .B0(N1017), .B1(n3785), .Y(n496) );
  NOR2XL U1904 ( .A(n3749), .B(\R[1][10] ), .Y(n3662) );
  NOR2XL U1905 ( .A(n3749), .B(\R[1][11] ), .Y(n3657) );
  NOR2XL U1906 ( .A(n3749), .B(\R[1][12] ), .Y(n3652) );
  AND4XL U1907 ( .A(n379), .B(n380), .C(n381), .D(n382), .Y(n134) );
  AND4XL U1908 ( .A(n373), .B(n374), .C(n375), .D(n376), .Y(n133) );
  NOR2XL U1909 ( .A(\R[3][10] ), .B(n3732), .Y(n3660) );
  NOR2XL U1910 ( .A(\R[3][11] ), .B(n3732), .Y(n3655) );
  NOR2XL U1911 ( .A(\R[3][12] ), .B(n3732), .Y(n3650) );
  MXI4XL U1912 ( .A(\R[28][10] ), .B(\R[29][10] ), .C(\R[30][10] ), .D(
        \R[31][10] ), .S0(n3718), .S1(n3743), .Y(n3339) );
  MXI4XL U1913 ( .A(\R[28][11] ), .B(\R[29][11] ), .C(\R[30][11] ), .D(
        \R[31][11] ), .S0(n3718), .S1(n3743), .Y(n3349) );
  MXI4XL U1914 ( .A(\R[28][12] ), .B(\R[29][12] ), .C(\R[30][12] ), .D(
        \R[31][12] ), .S0(n3718), .S1(n3743), .Y(n3359) );
  MXI4XL U1915 ( .A(\R[20][10] ), .B(\R[21][10] ), .C(\R[22][10] ), .D(
        \R[23][10] ), .S0(n3718), .S1(n3743), .Y(n3338) );
  MXI4XL U1916 ( .A(\R[4][10] ), .B(\R[5][10] ), .C(\R[6][10] ), .D(\R[7][10] ), .S0(n3718), .S1(n3743), .Y(n3343) );
  MXI4XL U1917 ( .A(\R[20][11] ), .B(\R[21][11] ), .C(\R[22][11] ), .D(
        \R[23][11] ), .S0(n3718), .S1(n3743), .Y(n3348) );
  MXI4XL U1918 ( .A(\R[4][11] ), .B(\R[5][11] ), .C(\R[6][11] ), .D(\R[7][11] ), .S0(n3718), .S1(n3743), .Y(n3353) );
  MXI4XL U1919 ( .A(\R[20][12] ), .B(\R[21][12] ), .C(\R[22][12] ), .D(
        \R[23][12] ), .S0(n3718), .S1(n3743), .Y(n3358) );
  MXI4XL U1920 ( .A(\R[4][12] ), .B(\R[5][12] ), .C(\R[6][12] ), .D(\R[7][12] ), .S0(n3718), .S1(n3743), .Y(n3363) );
  MXI4XL U1921 ( .A(\R[16][10] ), .B(\R[17][10] ), .C(\R[18][10] ), .D(
        \R[19][10] ), .S0(n3718), .S1(n3743), .Y(n3336) );
  MXI4XL U1922 ( .A(\R[16][11] ), .B(\R[17][11] ), .C(\R[18][11] ), .D(
        \R[19][11] ), .S0(n3718), .S1(n3743), .Y(n3346) );
  MXI4XL U1923 ( .A(\R[16][12] ), .B(\R[17][12] ), .C(\R[18][12] ), .D(
        \R[19][12] ), .S0(n3718), .S1(n3743), .Y(n3356) );
  MXI4XL U1924 ( .A(\R[8][10] ), .B(\R[9][10] ), .C(\R[10][10] ), .D(
        \R[11][10] ), .S0(n3718), .S1(n3743), .Y(n3342) );
  MXI4XL U1925 ( .A(\R[24][10] ), .B(\R[25][10] ), .C(\R[26][10] ), .D(
        \R[27][10] ), .S0(n3718), .S1(n3743), .Y(n3337) );
  MXI4XL U1926 ( .A(\R[8][11] ), .B(\R[9][11] ), .C(\R[10][11] ), .D(
        \R[11][11] ), .S0(n3718), .S1(n3743), .Y(n3352) );
  MXI4XL U1927 ( .A(\R[24][11] ), .B(\R[25][11] ), .C(\R[26][11] ), .D(
        \R[27][11] ), .S0(n3718), .S1(n3743), .Y(n3347) );
  MXI4XL U1928 ( .A(\R[8][12] ), .B(\R[9][12] ), .C(\R[10][12] ), .D(
        \R[11][12] ), .S0(n3718), .S1(n3743), .Y(n3362) );
  MXI4XL U1929 ( .A(\R[24][12] ), .B(\R[25][12] ), .C(\R[26][12] ), .D(
        \R[27][12] ), .S0(n3718), .S1(n3743), .Y(n3357) );
  NOR3X1 U1930 ( .A(instruction[26]), .B(instruction[27]), .C(instruction[25]), 
        .Y(n525) );
  NAND2X1 U1931 ( .A(n564), .B(n565), .Y(n465) );
  NOR3X1 U1932 ( .A(instruction[25]), .B(instruction[27]), .C(n4003), .Y(n551)
         );
  NOR2X1 U1933 ( .A(instruction[20]), .B(instruction[21]), .Y(n151) );
  NOR2X1 U1934 ( .A(n4007), .B(instruction[21]), .Y(n147) );
  CLKINVX1 U1935 ( .A(\seIM[31] ), .Y(n3972) );
  CLKINVX1 U1936 ( .A(N656), .Y(n3787) );
  CLKINVX1 U1937 ( .A(instruction[1]), .Y(n3974) );
  CLKINVX1 U1938 ( .A(instruction[2]), .Y(n3975) );
  CLKINVX1 U1939 ( .A(instruction[3]), .Y(n3976) );
  CLKINVX1 U1940 ( .A(instruction[4]), .Y(n3977) );
  CLKINVX1 U1941 ( .A(N52), .Y(n3981) );
  CLKINVX1 U1942 ( .A(N53), .Y(n3979) );
  CLKINVX1 U1943 ( .A(N54), .Y(n3978) );
  CLKINVX1 U1944 ( .A(N51), .Y(n3982) );
  CLKINVX1 U1945 ( .A(n3734), .Y(n3749) );
  CLKINVX1 U1946 ( .A(n3736), .Y(n3747) );
  CLKINVX1 U1947 ( .A(n3735), .Y(n3748) );
  CLKINVX1 U1948 ( .A(n3733), .Y(n3750) );
  CLKINVX1 U1949 ( .A(n3737), .Y(n3746) );
  INVX3 U1950 ( .A(n3740), .Y(n3743) );
  INVX3 U1951 ( .A(n3738), .Y(n3745) );
  INVX3 U1952 ( .A(n3739), .Y(n3744) );
  CLKINVX1 U1953 ( .A(n3741), .Y(n3742) );
  CLKINVX1 U1954 ( .A(n520), .Y(n4008) );
  CLKBUFX3 U1955 ( .A(n3725), .Y(n3719) );
  CLKBUFX3 U1956 ( .A(n3726), .Y(n3720) );
  BUFX4 U1957 ( .A(n3725), .Y(n3718) );
  BUFX4 U1958 ( .A(n3724), .Y(n3716) );
  BUFX4 U1959 ( .A(n3725), .Y(n3717) );
  CLKBUFX3 U1960 ( .A(n3726), .Y(n3721) );
  CLKBUFX3 U1961 ( .A(n3726), .Y(n3722) );
  CLKBUFX3 U1962 ( .A(n3724), .Y(n3715) );
  CLKBUFX3 U1963 ( .A(n3981), .Y(n3734) );
  CLKBUFX3 U1964 ( .A(n3981), .Y(n3735) );
  CLKBUFX3 U1965 ( .A(n3734), .Y(n3736) );
  CLKBUFX3 U1966 ( .A(n3735), .Y(n3737) );
  CLKBUFX3 U1967 ( .A(n3733), .Y(n3738) );
  CLKBUFX3 U1968 ( .A(n3736), .Y(n3739) );
  CLKBUFX3 U1969 ( .A(n3737), .Y(n3740) );
  CLKBUFX3 U1970 ( .A(n3981), .Y(n3733) );
  CLKBUFX3 U1971 ( .A(n3732), .Y(n3741) );
  CLKBUFX3 U1972 ( .A(n3736), .Y(n3732) );
  CLKBUFX3 U1973 ( .A(n3741), .Y(n3728) );
  CLKBUFX3 U1974 ( .A(n3741), .Y(n3729) );
  CLKBUFX3 U1975 ( .A(n3735), .Y(n3730) );
  CLKBUFX3 U1976 ( .A(n3737), .Y(n3731) );
  CLKBUFX3 U1977 ( .A(n3734), .Y(n3727) );
  CLKBUFX3 U1978 ( .A(n78), .Y(n3967) );
  CLKBUFX3 U1979 ( .A(n78), .Y(n3968) );
  CLKINVX1 U1980 ( .A(n3200), .Y(n3210) );
  CLKINVX1 U1981 ( .A(n3199), .Y(n3211) );
  CLKINVX1 U1982 ( .A(n3198), .Y(n3212) );
  CLKINVX1 U1983 ( .A(n3197), .Y(n3213) );
  CLKBUFX3 U1984 ( .A(n62), .Y(n3971) );
  NOR2X1 U1985 ( .A(n3210), .B(n3181), .Y(n3068) );
  NOR2X1 U1986 ( .A(n3210), .B(n3181), .Y(n3073) );
  NOR2X1 U1987 ( .A(n3210), .B(n3181), .Y(n3078) );
  NOR2X1 U1988 ( .A(n3211), .B(n3181), .Y(n3083) );
  NOR2X1 U1989 ( .A(n3211), .B(n3181), .Y(n3088) );
  NOR2X1 U1990 ( .A(n3211), .B(n3181), .Y(n3093) );
  NOR2X1 U1991 ( .A(n3211), .B(n3181), .Y(n3098) );
  NOR2X1 U1992 ( .A(n3211), .B(n3181), .Y(n3103) );
  NOR2X1 U1993 ( .A(n3211), .B(n3181), .Y(n3108) );
  NOR2X1 U1994 ( .A(n3212), .B(n3181), .Y(n3113) );
  NOR2X1 U1995 ( .A(n3212), .B(n3181), .Y(n3118) );
  NOR2X1 U1996 ( .A(n3212), .B(n3181), .Y(n3123) );
  INVX3 U1997 ( .A(n3202), .Y(n3209) );
  INVX3 U1998 ( .A(n3203), .Y(n3208) );
  INVX3 U1999 ( .A(n3204), .Y(n3207) );
  NOR2X1 U2000 ( .A(n3212), .B(n3182), .Y(n3018) );
  NOR2X1 U2001 ( .A(n3206), .B(n3182), .Y(n3023) );
  NOR2X1 U2002 ( .A(n3213), .B(n3182), .Y(n3028) );
  NOR2X1 U2003 ( .A(n3212), .B(n3182), .Y(n3033) );
  NOR2X1 U2004 ( .A(n3206), .B(n3182), .Y(n3038) );
  NOR2X1 U2005 ( .A(n3212), .B(n3182), .Y(n3043) );
  NOR2X1 U2006 ( .A(n3210), .B(n3182), .Y(n3048) );
  NOR2X1 U2007 ( .A(n3210), .B(n3182), .Y(n3053) );
  NOR2X1 U2008 ( .A(n3210), .B(n3182), .Y(n3058) );
  NOR2X1 U2009 ( .A(n3210), .B(n3182), .Y(n3063) );
  CLKBUFX3 U2010 ( .A(n78), .Y(n3969) );
  CLKINVX1 U2011 ( .A(n3205), .Y(n3206) );
  NOR2X1 U2012 ( .A(n3967), .B(n4024), .Y(address[0]) );
  NOR2X1 U2013 ( .A(n3967), .B(n4023), .Y(address[1]) );
  NOR2X1 U2014 ( .A(n3968), .B(n2683), .Y(address[2]) );
  NOR2X1 U2015 ( .A(n3968), .B(n2693), .Y(address[3]) );
  NOR2X1 U2016 ( .A(n3967), .B(n4017), .Y(address[10]) );
  NOR2X1 U2017 ( .A(n3967), .B(n4016), .Y(address[11]) );
  NOR2X1 U2018 ( .A(n3967), .B(n4015), .Y(address[12]) );
  NOR2X1 U2019 ( .A(n3967), .B(n2741), .Y(address[13]) );
  NOR2X1 U2020 ( .A(n3967), .B(n2750), .Y(address[14]) );
  NOR2X1 U2021 ( .A(n3967), .B(n4014), .Y(address[15]) );
  NOR2X1 U2022 ( .A(n3967), .B(n2713), .Y(address[16]) );
  NOR2X1 U2023 ( .A(n3967), .B(n2716), .Y(address[17]) );
  NOR2X1 U2024 ( .A(n3967), .B(n2710), .Y(address[18]) );
  NOR2X1 U2025 ( .A(n3967), .B(n4013), .Y(address[19]) );
  NOR2X1 U2026 ( .A(n3967), .B(n4012), .Y(address[20]) );
  NOR2X1 U2027 ( .A(n3968), .B(n2728), .Y(address[21]) );
  NOR2X1 U2028 ( .A(n3968), .B(n2707), .Y(address[22]) );
  NOR2X1 U2029 ( .A(n3968), .B(n2725), .Y(address[23]) );
  NOR2X1 U2030 ( .A(n3968), .B(n2699), .Y(address[24]) );
  NOR2X1 U2031 ( .A(n3968), .B(n4011), .Y(address[25]) );
  NOR2X1 U2032 ( .A(n3968), .B(n2704), .Y(address[26]) );
  NOR2X1 U2033 ( .A(n3968), .B(n4010), .Y(address[27]) );
  NOR2X1 U2034 ( .A(n3968), .B(n2696), .Y(address[28]) );
  NOR2X1 U2035 ( .A(n3968), .B(n2738), .Y(address[29]) );
  NOR2X1 U2036 ( .A(n3968), .B(n4009), .Y(address[30]) );
  NOR2X1 U2037 ( .A(n3968), .B(n2735), .Y(address[31]) );
  NOR2X1 U2038 ( .A(n3969), .B(n2686), .Y(address[4]) );
  NOR2X1 U2039 ( .A(n3969), .B(n4022), .Y(address[5]) );
  NOR2X1 U2040 ( .A(n3969), .B(n4021), .Y(address[6]) );
  NOR2X1 U2041 ( .A(n3969), .B(n4020), .Y(address[7]) );
  NOR2X1 U2042 ( .A(n3969), .B(n4019), .Y(address[8]) );
  NOR2X1 U2043 ( .A(n3969), .B(n4018), .Y(address[9]) );
  NAND2X1 U2044 ( .A(n526), .B(n527), .Y(n520) );
  NOR4X1 U2045 ( .A(n528), .B(n529), .C(n530), .D(n531), .Y(n527) );
  NOR4X1 U2046 ( .A(n532), .B(n533), .C(n534), .D(n535), .Y(n526) );
  NAND4X1 U2047 ( .A(n2693), .B(n2683), .C(n4023), .D(n4024), .Y(n528) );
  NAND4X1 U2048 ( .A(n4014), .B(n2750), .C(n2741), .D(n4015), .Y(n531) );
  NAND4X1 U2049 ( .A(n2735), .B(n4009), .C(n2738), .D(n2696), .Y(n535) );
  NAND4X1 U2050 ( .A(n4016), .B(n4017), .C(n4018), .D(n4019), .Y(n530) );
  NAND4X1 U2051 ( .A(n4010), .B(n2704), .C(n4011), .D(n2699), .Y(n534) );
  NAND4X1 U2052 ( .A(n4013), .B(n2710), .C(n2716), .D(n2713), .Y(n532) );
  NAND4X1 U2053 ( .A(n4020), .B(n4021), .C(n4022), .D(n2686), .Y(n529) );
  NAND4X1 U2054 ( .A(n2725), .B(n2707), .C(n2728), .D(n4012), .Y(n533) );
  CLKINVX1 U2055 ( .A(n3851), .Y(n3852) );
  CLKINVX1 U2056 ( .A(n3849), .Y(n3850) );
  CLKINVX1 U2057 ( .A(n3844), .Y(n3845) );
  CLKINVX1 U2058 ( .A(n3841), .Y(n3843) );
  CLKINVX1 U2059 ( .A(n3839), .Y(n3840) );
  CLKINVX1 U2060 ( .A(n3837), .Y(n3838) );
  CLKINVX1 U2061 ( .A(n3835), .Y(n3836) );
  CLKINVX1 U2062 ( .A(n3832), .Y(n3834) );
  CLKINVX1 U2063 ( .A(n3830), .Y(n3831) );
  CLKINVX1 U2064 ( .A(n3828), .Y(n3829) );
  CLKINVX1 U2065 ( .A(n3826), .Y(n3827) );
  CLKINVX1 U2066 ( .A(n3823), .Y(n3825) );
  CLKINVX1 U2067 ( .A(n3819), .Y(n3820) );
  CLKINVX1 U2068 ( .A(n3817), .Y(n3818) );
  CLKINVX1 U2069 ( .A(n3815), .Y(n3816) );
  CLKINVX1 U2070 ( .A(n3812), .Y(n3814) );
  CLKINVX1 U2071 ( .A(n3809), .Y(n3810) );
  CLKINVX1 U2072 ( .A(n3806), .Y(n3807) );
  CLKINVX1 U2073 ( .A(n3804), .Y(n3805) );
  CLKINVX1 U2074 ( .A(n3801), .Y(n3802) );
  CLKINVX1 U2075 ( .A(n3799), .Y(n3800) );
  CLKINVX1 U2076 ( .A(n3962), .Y(n3963) );
  CLKINVX1 U2077 ( .A(n3867), .Y(n3868) );
  CLKINVX1 U2078 ( .A(n3864), .Y(n3865) );
  CLKINVX1 U2079 ( .A(n3861), .Y(n3862) );
  CLKINVX1 U2080 ( .A(n3858), .Y(n3859) );
  CLKINVX1 U2081 ( .A(n3855), .Y(n3856) );
  CLKINVX1 U2082 ( .A(n3853), .Y(n3854) );
  CLKINVX1 U2083 ( .A(n3846), .Y(n3848) );
  CLKINVX1 U2084 ( .A(n3821), .Y(n3822) );
  CLKINVX1 U2085 ( .A(n3794), .Y(n3798) );
  CLKBUFX3 U2086 ( .A(n62), .Y(n3970) );
  CLKBUFX3 U2087 ( .A(n3770), .Y(n3768) );
  CLKBUFX3 U2088 ( .A(n3770), .Y(n3769) );
  CLKBUFX3 U2089 ( .A(n3765), .Y(n3761) );
  CLKBUFX3 U2090 ( .A(n3765), .Y(n3760) );
  CLKBUFX3 U2091 ( .A(n3766), .Y(n3764) );
  CLKBUFX3 U2092 ( .A(n3766), .Y(n3763) );
  CLKBUFX3 U2093 ( .A(n3766), .Y(n3762) );
  CLKBUFX3 U2094 ( .A(n3770), .Y(n3767) );
  CLKBUFX3 U2095 ( .A(n3723), .Y(n3726) );
  CLKBUFX3 U2096 ( .A(n3723), .Y(n3725) );
  CLKBUFX3 U2097 ( .A(n3757), .Y(n3753) );
  CLKBUFX3 U2098 ( .A(n3757), .Y(n3752) );
  CLKBUFX3 U2099 ( .A(n3758), .Y(n3756) );
  CLKBUFX3 U2100 ( .A(n3758), .Y(n3755) );
  CLKBUFX3 U2101 ( .A(n3758), .Y(n3754) );
  CLKBUFX3 U2102 ( .A(n3723), .Y(n3724) );
  CLKBUFX3 U2103 ( .A(n3765), .Y(n3759) );
  CLKBUFX3 U2104 ( .A(n3757), .Y(n3751) );
  AOI222XL U2105 ( .A0(N431), .A1(n250), .B0(N623), .B1(n248), .C0(N463), .C1(
        n246), .Y(n313) );
  AOI222XL U2106 ( .A0(N430), .A1(n3779), .B0(N622), .B1(n3780), .C0(N462), 
        .C1(n246), .Y(n327) );
  AOI222XL U2107 ( .A0(N429), .A1(n250), .B0(N621), .B1(n248), .C0(N461), .C1(
        n246), .Y(n333) );
  AOI222XL U2108 ( .A0(N428), .A1(n3779), .B0(N620), .B1(n3780), .C0(N460), 
        .C1(n246), .Y(n339) );
  AOI222XL U2109 ( .A0(N427), .A1(n250), .B0(N619), .B1(n248), .C0(N459), .C1(
        n246), .Y(n345) );
  CLKBUFX3 U2110 ( .A(n3188), .Y(n3182) );
  BUFX4 U2111 ( .A(n3186), .Y(n3178) );
  BUFX4 U2112 ( .A(n3187), .Y(n3180) );
  BUFX4 U2113 ( .A(n3187), .Y(n3179) );
  CLKBUFX3 U2114 ( .A(n3188), .Y(n3183) );
  CLKBUFX3 U2115 ( .A(n3188), .Y(n3184) );
  NAND2BX1 U2116 ( .AN(n111), .B(n4045), .Y(n62) );
  CLKBUFX3 U2117 ( .A(n3186), .Y(n3177) );
  AND2X2 U2118 ( .A(MR), .B(n3971), .Y(n78) );
  CLKBUFX3 U2119 ( .A(n3190), .Y(n3201) );
  CLKBUFX3 U2120 ( .A(n3190), .Y(n3200) );
  CLKBUFX3 U2121 ( .A(n3200), .Y(n3199) );
  CLKBUFX3 U2122 ( .A(n3190), .Y(n3198) );
  CLKBUFX3 U2123 ( .A(n3201), .Y(n3197) );
  CLKBUFX3 U2124 ( .A(n3189), .Y(n3205) );
  CLKBUFX3 U2125 ( .A(n3190), .Y(n3202) );
  CLKBUFX3 U2126 ( .A(n3189), .Y(n3203) );
  CLKBUFX3 U2127 ( .A(n3189), .Y(n3204) );
  CLKBUFX3 U2128 ( .A(n3197), .Y(n3192) );
  CLKBUFX3 U2129 ( .A(n3198), .Y(n3193) );
  CLKBUFX3 U2130 ( .A(n3195), .Y(n3194) );
  CLKBUFX3 U2131 ( .A(n3205), .Y(n3195) );
  CLKBUFX3 U2132 ( .A(n3197), .Y(n3196) );
  CLKBUFX3 U2133 ( .A(n3197), .Y(n3191) );
  INVX1 U2134 ( .A(n2648), .Y(n4012) );
  INVX1 U2135 ( .A(n2651), .Y(n4010) );
  INVX1 U2136 ( .A(n2649), .Y(n4013) );
  INVX1 U2137 ( .A(n2653), .Y(n4014) );
  INVX1 U2138 ( .A(n2670), .Y(n4024) );
  INVX1 U2139 ( .A(n2650), .Y(n4011) );
  INVX1 U2140 ( .A(n2652), .Y(n4009) );
  CLKINVX1 U2141 ( .A(n2676), .Y(n4016) );
  CLKINVX1 U2142 ( .A(n2677), .Y(n4015) );
  CLKINVX1 U2143 ( .A(n2675), .Y(n4019) );
  CLKINVX1 U2144 ( .A(n2674), .Y(n4018) );
  CLKINVX1 U2145 ( .A(n2655), .Y(n4022) );
  CLKINVX1 U2146 ( .A(n2673), .Y(n4017) );
  CLKINVX1 U2147 ( .A(n2671), .Y(n4020) );
  CLKINVX1 U2148 ( .A(n2672), .Y(n4021) );
  AOI222XL U2149 ( .A0(N426), .A1(n3779), .B0(N618), .B1(n3780), .C0(N458), 
        .C1(n3774), .Y(n351) );
  AOI222XL U2150 ( .A0(N425), .A1(n250), .B0(N617), .B1(n248), .C0(N457), .C1(
        n246), .Y(n357) );
  AOI222XL U2151 ( .A0(N424), .A1(n3779), .B0(N616), .B1(n3780), .C0(N456), 
        .C1(n3774), .Y(n363) );
  AOI222XL U2152 ( .A0(N423), .A1(n250), .B0(N615), .B1(n248), .C0(N455), .C1(
        n246), .Y(n369) );
  AOI222XL U2153 ( .A0(N422), .A1(n3779), .B0(N614), .B1(n3780), .C0(N454), 
        .C1(n3774), .Y(n375) );
  AOI222XL U2154 ( .A0(N421), .A1(n250), .B0(N613), .B1(n248), .C0(N453), .C1(
        n246), .Y(n381) );
  AOI222XL U2155 ( .A0(N447), .A1(n3774), .B0(N671), .B1(n3781), .C0(N607), 
        .C1(n248), .Y(n425) );
  AOI222XL U2156 ( .A0(N420), .A1(n3779), .B0(N612), .B1(n3780), .C0(N452), 
        .C1(n3774), .Y(n395) );
  AOI222XL U2157 ( .A0(N419), .A1(n250), .B0(N611), .B1(n248), .C0(N451), .C1(
        n246), .Y(n401) );
  AOI222XL U2158 ( .A0(N418), .A1(n3779), .B0(N610), .B1(n3780), .C0(N450), 
        .C1(n3774), .Y(n407) );
  AOI222XL U2159 ( .A0(N417), .A1(n250), .B0(N609), .B1(n248), .C0(N449), .C1(
        n246), .Y(n413) );
  AOI222XL U2160 ( .A0(N416), .A1(n3779), .B0(N608), .B1(n3780), .C0(N448), 
        .C1(n3774), .Y(n419) );
  CLKBUFX3 U2161 ( .A(n121), .Y(n3944) );
  CLKBUFX3 U2162 ( .A(n121), .Y(n3945) );
  AOI222XL U2163 ( .A0(N446), .A1(n246), .B0(N670), .B1(n247), .C0(N606), .C1(
        n3780), .Y(n433) );
  AOI222XL U2164 ( .A0(N445), .A1(n3774), .B0(N669), .B1(n3781), .C0(N605), 
        .C1(n248), .Y(n441) );
  AOI222XL U2165 ( .A0(N444), .A1(n246), .B0(N668), .B1(n247), .C0(N604), .C1(
        n3780), .Y(n449) );
  AOI222XL U2166 ( .A0(N443), .A1(n3774), .B0(N667), .B1(n3781), .C0(N603), 
        .C1(n248), .Y(n457) );
  CLKBUFX3 U2167 ( .A(n121), .Y(n3946) );
  CLKBUFX3 U2168 ( .A(n120), .Y(n3947) );
  CLKBUFX3 U2169 ( .A(n124), .Y(n3935) );
  CLKBUFX3 U2170 ( .A(n135), .Y(n3902) );
  CLKBUFX3 U2171 ( .A(n120), .Y(n3948) );
  CLKBUFX3 U2172 ( .A(n124), .Y(n3936) );
  CLKBUFX3 U2173 ( .A(n135), .Y(n3903) );
  CLKBUFX3 U2174 ( .A(n3993), .Y(n3784) );
  CLKBUFX3 U2175 ( .A(n3993), .Y(n3785) );
  CLKBUFX3 U2176 ( .A(n3993), .Y(n3786) );
  CLKBUFX3 U2177 ( .A(n120), .Y(n3949) );
  CLKBUFX3 U2178 ( .A(n124), .Y(n3937) );
  CLKBUFX3 U2179 ( .A(n135), .Y(n3904) );
  CLKBUFX3 U2180 ( .A(n2654), .Y(n3973) );
  CLKBUFX3 U2181 ( .A(n228), .Y(n3796) );
  CLKBUFX3 U2182 ( .A(n228), .Y(n3795) );
  CLKBUFX3 U2183 ( .A(n228), .Y(n3794) );
  CLKBUFX3 U2184 ( .A(n228), .Y(n3797) );
  CLKBUFX3 U2185 ( .A(n114), .Y(n3962) );
  CLKBUFX3 U2186 ( .A(n149), .Y(n3867) );
  CLKBUFX3 U2187 ( .A(n175), .Y(n3844) );
  CLKBUFX3 U2188 ( .A(n186), .Y(n3835) );
  CLKBUFX3 U2189 ( .A(n196), .Y(n3826) );
  CLKBUFX3 U2190 ( .A(n209), .Y(n3815) );
  CLKBUFX3 U2191 ( .A(n219), .Y(n3804) );
  CLKBUFX3 U2192 ( .A(n201), .Y(n3821) );
  CLKBUFX3 U2193 ( .A(n177), .Y(n3841) );
  CLKBUFX3 U2194 ( .A(n188), .Y(n3832) );
  CLKBUFX3 U2195 ( .A(n198), .Y(n3823) );
  CLKBUFX3 U2196 ( .A(n211), .Y(n3812) );
  CLKBUFX3 U2197 ( .A(n225), .Y(n3799) );
  CLKBUFX3 U2198 ( .A(n168), .Y(n3851) );
  CLKBUFX3 U2199 ( .A(n171), .Y(n3849) );
  CLKBUFX3 U2200 ( .A(n181), .Y(n3839) );
  CLKBUFX3 U2201 ( .A(n184), .Y(n3837) );
  CLKBUFX3 U2202 ( .A(n191), .Y(n3830) );
  CLKBUFX3 U2203 ( .A(n194), .Y(n3828) );
  CLKBUFX3 U2204 ( .A(n204), .Y(n3819) );
  CLKBUFX3 U2205 ( .A(n207), .Y(n3817) );
  CLKBUFX3 U2206 ( .A(n165), .Y(n3853) );
  CLKBUFX3 U2207 ( .A(n173), .Y(n3846) );
  CLKBUFX3 U2208 ( .A(n480), .Y(n3788) );
  CLKBUFX3 U2209 ( .A(n480), .Y(n3789) );
  CLKBUFX3 U2210 ( .A(n177), .Y(n3842) );
  CLKBUFX3 U2211 ( .A(n188), .Y(n3833) );
  CLKBUFX3 U2212 ( .A(n198), .Y(n3824) );
  CLKBUFX3 U2213 ( .A(n211), .Y(n3813) );
  CLKINVX1 U2214 ( .A(n3809), .Y(n3811) );
  CLKBUFX3 U2215 ( .A(n214), .Y(n3809) );
  CLKINVX1 U2216 ( .A(n3806), .Y(n3808) );
  CLKBUFX3 U2217 ( .A(n217), .Y(n3806) );
  CLKINVX1 U2218 ( .A(n3801), .Y(n3803) );
  CLKBUFX3 U2219 ( .A(n222), .Y(n3801) );
  CLKINVX1 U2220 ( .A(n3864), .Y(n3866) );
  CLKBUFX3 U2221 ( .A(n152), .Y(n3864) );
  CLKINVX1 U2222 ( .A(n3861), .Y(n3863) );
  CLKBUFX3 U2223 ( .A(n156), .Y(n3861) );
  CLKINVX1 U2224 ( .A(n3858), .Y(n3860) );
  CLKBUFX3 U2225 ( .A(n159), .Y(n3858) );
  CLKINVX1 U2226 ( .A(n3855), .Y(n3857) );
  CLKBUFX3 U2227 ( .A(n161), .Y(n3855) );
  CLKBUFX3 U2228 ( .A(n173), .Y(n3847) );
  CLKBUFX3 U2229 ( .A(n480), .Y(n3790) );
  OAI221XL U2230 ( .A0(n2735), .A1(n3773), .B0(N190), .B1(n3792), .C0(n3996), 
        .Y(n308) );
  OAI221XL U2231 ( .A0(n4009), .A1(n238), .B0(n2652), .B1(n3792), .C0(n3996), 
        .Y(n316) );
  OAI221XL U2232 ( .A0(n2738), .A1(n238), .B0(N192), .B1(n3792), .C0(n3996), 
        .Y(n330) );
  OAI221XL U2233 ( .A0(n2696), .A1(n3773), .B0(N193), .B1(n3792), .C0(n3996), 
        .Y(n336) );
  OAI221XL U2234 ( .A0(n4010), .A1(n238), .B0(n2651), .B1(n3792), .C0(n3996), 
        .Y(n342) );
  OAI221XL U2235 ( .A0(n2704), .A1(n3773), .B0(N195), .B1(n3792), .C0(n3996), 
        .Y(n348) );
  OAI221XL U2236 ( .A0(n4011), .A1(n238), .B0(n2650), .B1(n3792), .C0(n3996), 
        .Y(n354) );
  OAI221XL U2237 ( .A0(n2699), .A1(n3773), .B0(N197), .B1(n3792), .C0(n3996), 
        .Y(n360) );
  OAI221XL U2238 ( .A0(n2725), .A1(n238), .B0(N198), .B1(n3792), .C0(n3996), 
        .Y(n366) );
  OAI221XL U2239 ( .A0(n2707), .A1(n3773), .B0(N199), .B1(n3792), .C0(n3996), 
        .Y(n372) );
  OAI221XL U2240 ( .A0(n2728), .A1(n238), .B0(N200), .B1(n3792), .C0(n3996), 
        .Y(n378) );
  OAI221XL U2241 ( .A0(n4012), .A1(n3773), .B0(n2648), .B1(n3792), .C0(n3996), 
        .Y(n384) );
  OAI221XL U2242 ( .A0(n4013), .A1(n3773), .B0(n2649), .B1(n3792), .C0(n3996), 
        .Y(n398) );
  OAI221XL U2243 ( .A0(n2710), .A1(n238), .B0(N203), .B1(n3792), .C0(n3996), 
        .Y(n404) );
  OAI221XL U2244 ( .A0(n2716), .A1(n3773), .B0(N204), .B1(n3792), .C0(n3996), 
        .Y(n410) );
  OAI221XL U2245 ( .A0(n2713), .A1(n238), .B0(N205), .B1(n3792), .C0(n3996), 
        .Y(n416) );
  OAI221XL U2246 ( .A0(n4014), .A1(n3773), .B0(n2653), .B1(n3792), .C0(n3996), 
        .Y(n422) );
  NOR4BBX1 U2247 ( .AN(n3773), .BN(n3792), .C(n3774), .D(n242), .Y(n547) );
  CLKINVX1 U2248 ( .A(n462), .Y(n3996) );
  CLKBUFX3 U2249 ( .A(n239), .Y(n3792) );
  CLKBUFX3 U2250 ( .A(n239), .Y(n3791) );
  CLKINVX1 U2251 ( .A(n244), .Y(n3998) );
  NOR2X1 U2252 ( .A(n3970), .B(n4039), .Y(datain[0]) );
  NOR2X1 U2253 ( .A(n3970), .B(n4037), .Y(datain[2]) );
  NOR2X1 U2254 ( .A(n3970), .B(n4036), .Y(datain[3]) );
  NOR2X1 U2255 ( .A(n3970), .B(n4035), .Y(datain[4]) );
  NOR2X1 U2256 ( .A(n3970), .B(n4034), .Y(datain[5]) );
  NOR2X1 U2257 ( .A(n3970), .B(n4033), .Y(datain[6]) );
  NOR2X1 U2258 ( .A(n3970), .B(n4032), .Y(datain[7]) );
  NOR2X1 U2259 ( .A(n3970), .B(n4031), .Y(datain[8]) );
  NOR2X1 U2260 ( .A(n3970), .B(n4030), .Y(datain[9]) );
  NOR2X1 U2261 ( .A(n3970), .B(n4029), .Y(datain[10]) );
  NOR2X1 U2262 ( .A(n3970), .B(n4028), .Y(datain[11]) );
  NOR2X1 U2263 ( .A(n3970), .B(n4027), .Y(datain[12]) );
  NOR2X1 U2264 ( .A(n3970), .B(n4026), .Y(datain[13]) );
  CLKBUFX3 U2265 ( .A(\seIM[31] ), .Y(n3770) );
  NOR2X1 U2266 ( .A(n3971), .B(n4038), .Y(datain[1]) );
  NOR2X1 U2267 ( .A(n3971), .B(n4025), .Y(datain[14]) );
  CLKBUFX3 U2268 ( .A(N54), .Y(n3765) );
  CLKBUFX3 U2269 ( .A(N53), .Y(n3757) );
  CLKBUFX3 U2270 ( .A(N54), .Y(n3766) );
  CLKBUFX3 U2271 ( .A(N53), .Y(n3758) );
  CLKBUFX3 U2272 ( .A(N51), .Y(n3723) );
  CLKBUFX3 U2273 ( .A(n239), .Y(n3793) );
  CLKBUFX3 U2274 ( .A(n122), .Y(n3941) );
  CLKBUFX3 U2275 ( .A(n122), .Y(n3942) );
  MX4X1 U2276 ( .A(n2773), .B(n2774), .C(n2775), .D(n2776), .S0(n3223), .S1(
        n3215), .Y(n2679) );
  NAND2X1 U2277 ( .A(n3171), .B(n3170), .Y(n2773) );
  NOR2X1 U2278 ( .A(n3169), .B(n3168), .Y(n3171) );
  MXI2X1 U2279 ( .A(n1532), .B(n3167), .S0(n3184), .Y(n3170) );
  NOR2X1 U2280 ( .A(n3213), .B(n3181), .Y(n3168) );
  MX4X1 U2281 ( .A(n2801), .B(n2802), .C(n2803), .D(n2804), .S0(n3224), .S1(
        n3216), .Y(n2690) );
  CLKBUFX3 U2282 ( .A(n123), .Y(n3938) );
  CLKBUFX3 U2283 ( .A(n125), .Y(n3932) );
  CLKBUFX3 U2284 ( .A(n126), .Y(n3929) );
  CLKBUFX3 U2285 ( .A(n127), .Y(n3926) );
  CLKBUFX3 U2286 ( .A(n128), .Y(n3923) );
  CLKBUFX3 U2287 ( .A(n123), .Y(n3939) );
  CLKBUFX3 U2288 ( .A(n125), .Y(n3933) );
  CLKBUFX3 U2289 ( .A(n126), .Y(n3930) );
  CLKBUFX3 U2290 ( .A(n127), .Y(n3927) );
  CLKBUFX3 U2291 ( .A(n128), .Y(n3924) );
  MX4X1 U2292 ( .A(n2813), .B(n2814), .C(n2815), .D(n2816), .S0(n3224), .S1(
        n3216), .Y(n2691) );
  MX4X1 U2293 ( .A(n2809), .B(n2810), .C(n2811), .D(n2812), .S0(n3224), .S1(
        n3216), .Y(n2692) );
  CLKBUFX3 U2294 ( .A(n123), .Y(n3940) );
  CLKBUFX3 U2295 ( .A(n125), .Y(n3934) );
  CLKBUFX3 U2296 ( .A(n126), .Y(n3931) );
  NAND2X1 U2297 ( .A(n3176), .B(n3175), .Y(n2765) );
  NOR2X1 U2298 ( .A(n3174), .B(n3173), .Y(n3176) );
  MXI2X1 U2299 ( .A(n1533), .B(n3172), .S0(n3184), .Y(n3175) );
  NOR2X1 U2300 ( .A(n3213), .B(n3181), .Y(n3173) );
  NAND2X1 U2301 ( .A(n3146), .B(n3145), .Y(n2813) );
  NOR2X1 U2302 ( .A(n3144), .B(n3143), .Y(n3146) );
  MXI2X1 U2303 ( .A(n1527), .B(n3142), .S0(n3184), .Y(n3145) );
  NOR2X1 U2304 ( .A(n3212), .B(n3181), .Y(n3143) );
  NAND2X1 U2305 ( .A(n3151), .B(n3150), .Y(n2805) );
  NOR2X1 U2306 ( .A(n3149), .B(n3148), .Y(n3151) );
  MXI2X1 U2307 ( .A(n1528), .B(n3147), .S0(n3184), .Y(n3150) );
  NOR2X1 U2308 ( .A(n3213), .B(n3181), .Y(n3148) );
  NAND2X1 U2309 ( .A(n3689), .B(n3688), .Y(n3291) );
  NOR2X1 U2310 ( .A(n3687), .B(n3686), .Y(n3689) );
  MXI2X1 U2311 ( .A(n1528), .B(n3685), .S0(n3722), .Y(n3688) );
  NOR2X1 U2312 ( .A(n3750), .B(n3719), .Y(n3686) );
  NAND2X1 U2313 ( .A(n3156), .B(n3155), .Y(n2797) );
  NOR2X1 U2314 ( .A(n3154), .B(n3153), .Y(n3156) );
  MXI2X1 U2315 ( .A(n1529), .B(n3152), .S0(n3184), .Y(n3155) );
  NOR2X1 U2316 ( .A(n3213), .B(n3181), .Y(n3153) );
  NAND2X1 U2317 ( .A(n3694), .B(n3693), .Y(n3281) );
  NOR2X1 U2318 ( .A(n3692), .B(n3691), .Y(n3694) );
  MXI2X1 U2319 ( .A(n1529), .B(n3690), .S0(n3722), .Y(n3693) );
  NOR2X1 U2320 ( .A(n3750), .B(n3719), .Y(n3691) );
  NAND2X1 U2321 ( .A(n3161), .B(n3160), .Y(n2789) );
  NOR2X1 U2322 ( .A(n3159), .B(n3158), .Y(n3161) );
  MXI2X1 U2323 ( .A(n1530), .B(n3157), .S0(n3184), .Y(n3160) );
  NOR2X1 U2324 ( .A(n3213), .B(n3181), .Y(n3158) );
  NAND2X1 U2325 ( .A(n3699), .B(n3698), .Y(n3271) );
  NOR2X1 U2326 ( .A(n3697), .B(n3696), .Y(n3699) );
  MXI2X1 U2327 ( .A(n1530), .B(n3695), .S0(n3722), .Y(n3698) );
  NOR2X1 U2328 ( .A(n3750), .B(n3719), .Y(n3696) );
  NAND2X1 U2329 ( .A(n3166), .B(n3165), .Y(n2781) );
  NOR2X1 U2330 ( .A(n3164), .B(n3163), .Y(n3166) );
  MXI2X1 U2331 ( .A(n1531), .B(n3162), .S0(n3184), .Y(n3165) );
  NOR2X1 U2332 ( .A(n3213), .B(n3181), .Y(n3163) );
  NAND2X1 U2333 ( .A(n3704), .B(n3703), .Y(n3261) );
  NOR2X1 U2334 ( .A(n3702), .B(n3701), .Y(n3704) );
  MXI2X1 U2335 ( .A(n1531), .B(n3700), .S0(n3722), .Y(n3703) );
  NOR2X1 U2336 ( .A(n3750), .B(n3719), .Y(n3701) );
  NAND2X1 U2337 ( .A(n3709), .B(n3708), .Y(n3251) );
  NOR2X1 U2338 ( .A(n3707), .B(n3706), .Y(n3709) );
  MXI2X1 U2339 ( .A(n1532), .B(n3705), .S0(n3722), .Y(n3708) );
  NOR2X1 U2340 ( .A(n3750), .B(n3719), .Y(n3706) );
  NAND2X1 U2341 ( .A(n3714), .B(n3713), .Y(n3241) );
  NOR2X1 U2342 ( .A(n3712), .B(n3711), .Y(n3714) );
  MXI2X1 U2343 ( .A(n1533), .B(n3710), .S0(n3722), .Y(n3713) );
  NOR2X1 U2344 ( .A(n3750), .B(n3719), .Y(n3711) );
  AND2X2 U2345 ( .A(n543), .B(n3994), .Y(n524) );
  CLKMX2X2 U2346 ( .A(n2697), .B(n2698), .S0(n3233), .Y(n2696) );
  CLKINVX1 U2347 ( .A(n2696), .Y(N193) );
  MX4X1 U2348 ( .A(n2989), .B(n2990), .C(n2991), .D(n2992), .S0(n3228), .S1(
        n3220), .Y(n2697) );
  MX4X1 U2349 ( .A(n2985), .B(n2986), .C(n2987), .D(n2988), .S0(n3228), .S1(
        n3220), .Y(n2698) );
  NAND2X1 U2350 ( .A(n524), .B(n525), .Y(n111) );
  CLKMX2X2 U2351 ( .A(n2700), .B(n2701), .S0(n3233), .Y(n2699) );
  CLKINVX1 U2352 ( .A(n2699), .Y(N197) );
  MX4X1 U2353 ( .A(n2957), .B(n2958), .C(n2959), .D(n2960), .S0(n3227), .S1(
        n3219), .Y(n2700) );
  MX4X1 U2354 ( .A(n2953), .B(n2954), .C(n2955), .D(n2956), .S0(n3227), .S1(
        n3219), .Y(n2701) );
  MX4X1 U2355 ( .A(n2925), .B(n2926), .C(n2927), .D(n2928), .S0(n3227), .S1(
        n3219), .Y(n2702) );
  MX4X1 U2356 ( .A(n2921), .B(n2922), .C(n2923), .D(n2924), .S0(n3227), .S1(
        n3219), .Y(n2703) );
  CLKMX2X2 U2357 ( .A(n2705), .B(n2706), .S0(n3233), .Y(n2704) );
  CLKINVX1 U2358 ( .A(n2704), .Y(N195) );
  MX4X1 U2359 ( .A(n2973), .B(n2974), .C(n2975), .D(n2976), .S0(n3228), .S1(
        n3220), .Y(n2705) );
  MX4X1 U2360 ( .A(n2969), .B(n2970), .C(n2971), .D(n2972), .S0(n3228), .S1(
        n3220), .Y(n2706) );
  CLKMX2X2 U2361 ( .A(n2708), .B(n2709), .S0(n3233), .Y(n2707) );
  MX4X1 U2362 ( .A(n2941), .B(n2942), .C(n2943), .D(n2944), .S0(n3227), .S1(
        n3219), .Y(n2708) );
  MX4X1 U2363 ( .A(n2937), .B(n2938), .C(n2939), .D(n2940), .S0(n3227), .S1(
        n3219), .Y(n2709) );
  CLKMX2X2 U2364 ( .A(n2711), .B(n2712), .S0(n3232), .Y(n2710) );
  CLKINVX1 U2365 ( .A(n2710), .Y(N203) );
  MX4X1 U2366 ( .A(n2909), .B(n2910), .C(n2911), .D(n2912), .S0(n3226), .S1(
        n3218), .Y(n2711) );
  MX4X1 U2367 ( .A(n2905), .B(n2906), .C(n2907), .D(n2908), .S0(n3226), .S1(
        n3218), .Y(n2712) );
  CLKMX2X2 U2368 ( .A(n2714), .B(n2715), .S0(n3232), .Y(n2713) );
  CLKINVX1 U2369 ( .A(n2713), .Y(N205) );
  MX4X1 U2370 ( .A(n2893), .B(n2894), .C(n2895), .D(n2896), .S0(n3226), .S1(
        n3218), .Y(n2714) );
  MX4X1 U2371 ( .A(n2889), .B(n2890), .C(n2891), .D(n2892), .S0(n3226), .S1(
        n3218), .Y(n2715) );
  CLKMX2X2 U2372 ( .A(n2717), .B(n2718), .S0(n3232), .Y(n2716) );
  CLKINVX1 U2373 ( .A(n2716), .Y(N204) );
  MX4X1 U2374 ( .A(n2901), .B(n2902), .C(n2903), .D(n2904), .S0(n3226), .S1(
        n3218), .Y(n2717) );
  MX4X1 U2375 ( .A(n2897), .B(n2898), .C(n2899), .D(n2900), .S0(n3226), .S1(
        n3218), .Y(n2718) );
  MX4X1 U2376 ( .A(n3005), .B(n3006), .C(n3007), .D(n3008), .S0(n3228), .S1(
        n3220), .Y(n2719) );
  MX4X1 U2377 ( .A(n3001), .B(n3002), .C(n3003), .D(n3004), .S0(n3228), .S1(
        n3220), .Y(n2720) );
  MX4X1 U2378 ( .A(n2981), .B(n2982), .C(n2983), .D(n2984), .S0(n3228), .S1(
        n3220), .Y(n2721) );
  MX4X1 U2379 ( .A(n2977), .B(n2978), .C(n2979), .D(n2980), .S0(n3228), .S1(
        n3220), .Y(n2722) );
  MX4X1 U2380 ( .A(n2965), .B(n2966), .C(n2967), .D(n2968), .S0(n3227), .S1(
        n3219), .Y(n2723) );
  MX4X1 U2381 ( .A(n2961), .B(n2962), .C(n2963), .D(n2964), .S0(n3227), .S1(
        n3219), .Y(n2724) );
  CLKMX2X2 U2382 ( .A(n2726), .B(n2727), .S0(n3233), .Y(n2725) );
  MX4X1 U2383 ( .A(n2949), .B(n2950), .C(n2951), .D(n2952), .S0(n3227), .S1(
        n3219), .Y(n2726) );
  MX4X1 U2384 ( .A(n2945), .B(n2946), .C(n2947), .D(n2948), .S0(n3227), .S1(
        n3219), .Y(n2727) );
  CLKMX2X2 U2385 ( .A(n2729), .B(n2730), .S0(n3233), .Y(n2728) );
  CLKINVX1 U2386 ( .A(n2728), .Y(N200) );
  MX4X1 U2387 ( .A(n2933), .B(n2934), .C(n2935), .D(n2936), .S0(n3227), .S1(
        n3219), .Y(n2729) );
  MX4X1 U2388 ( .A(n2929), .B(n2930), .C(n2931), .D(n2932), .S0(n3227), .S1(
        n3219), .Y(n2730) );
  MX4X1 U2389 ( .A(n2917), .B(n2918), .C(n2919), .D(n2920), .S0(n3226), .S1(
        n3218), .Y(n2731) );
  MX4X1 U2390 ( .A(n2913), .B(n2914), .C(n2915), .D(n2916), .S0(n3226), .S1(
        n3218), .Y(n2732) );
  MX4X1 U2391 ( .A(n2885), .B(n2886), .C(n2887), .D(n2888), .S0(n3226), .S1(
        n3218), .Y(n2733) );
  MX4X1 U2392 ( .A(n2881), .B(n2882), .C(n2883), .D(n2884), .S0(n3226), .S1(
        n3218), .Y(n2734) );
  CLKMX2X2 U2393 ( .A(n2736), .B(n2737), .S0(n3233), .Y(n2735) );
  CLKINVX1 U2394 ( .A(n2735), .Y(N190) );
  MX4X1 U2395 ( .A(n3013), .B(n3014), .C(n3015), .D(n3016), .S0(n3228), .S1(
        n3220), .Y(n2736) );
  MX4X1 U2396 ( .A(n3009), .B(n3010), .C(n3011), .D(n3012), .S0(n3228), .S1(
        n3220), .Y(n2737) );
  CLKMX2X2 U2397 ( .A(n2739), .B(n2740), .S0(n3233), .Y(n2738) );
  CLKINVX1 U2398 ( .A(n2738), .Y(N192) );
  MX4X1 U2399 ( .A(n2997), .B(n2998), .C(n2999), .D(n3000), .S0(n3228), .S1(
        n3220), .Y(n2739) );
  MX4X1 U2400 ( .A(n2993), .B(n2994), .C(n2995), .D(n2996), .S0(n3228), .S1(
        n3220), .Y(n2740) );
  CLKMX2X2 U2401 ( .A(n2742), .B(n2743), .S0(n3232), .Y(n2741) );
  CLKINVX1 U2402 ( .A(n2741), .Y(N208) );
  MX4X1 U2403 ( .A(n2869), .B(n2870), .C(n2871), .D(n2872), .S0(n3225), .S1(
        n3217), .Y(n2742) );
  MX4X1 U2404 ( .A(n2865), .B(n2866), .C(n2867), .D(n2868), .S0(n3225), .S1(
        n3217), .Y(n2743) );
  MX4X1 U2405 ( .A(n2861), .B(n2862), .C(n2863), .D(n2864), .S0(n3225), .S1(
        n3217), .Y(n2744) );
  MX4X1 U2406 ( .A(n2857), .B(n2858), .C(n2859), .D(n2860), .S0(n3225), .S1(
        n3217), .Y(n2745) );
  MX4X1 U2407 ( .A(n2853), .B(n2854), .C(n2855), .D(n2856), .S0(n3225), .S1(
        n3217), .Y(n2746) );
  MX4X1 U2408 ( .A(n2849), .B(n2850), .C(n2851), .D(n2852), .S0(n3225), .S1(
        n3217), .Y(n2747) );
  MX4X1 U2409 ( .A(n2845), .B(n2846), .C(n2847), .D(n2848), .S0(n3225), .S1(
        n3217), .Y(n2748) );
  AND2X2 U2410 ( .A(n539), .B(n3999), .Y(n3771) );
  CLKBUFX3 U2411 ( .A(n129), .Y(n3920) );
  CLKBUFX3 U2412 ( .A(n133), .Y(n3908) );
  CLKBUFX3 U2413 ( .A(n134), .Y(n3905) );
  CLKBUFX3 U2414 ( .A(n129), .Y(n3921) );
  CLKBUFX3 U2415 ( .A(n133), .Y(n3909) );
  CLKBUFX3 U2416 ( .A(n134), .Y(n3906) );
  CLKMX2X2 U2417 ( .A(n2751), .B(n2752), .S0(n3232), .Y(n2750) );
  MX4X1 U2418 ( .A(n2877), .B(n2878), .C(n2879), .D(n2880), .S0(n3226), .S1(
        n3218), .Y(n2751) );
  MX4X1 U2419 ( .A(n2873), .B(n2874), .C(n2875), .D(n2876), .S0(n3226), .S1(
        n3218), .Y(n2752) );
  CLKBUFX3 U2420 ( .A(n3230), .Y(n3228) );
  CLKBUFX3 U2421 ( .A(n3230), .Y(n3227) );
  CLKBUFX3 U2422 ( .A(n3230), .Y(n3226) );
  CLKBUFX3 U2423 ( .A(n3229), .Y(n3225) );
  CLKBUFX3 U2424 ( .A(n3229), .Y(n3224) );
  MX4X1 U2425 ( .A(n2837), .B(n2838), .C(n2839), .D(n2840), .S0(n3225), .S1(
        n3217), .Y(n2753) );
  MX4X1 U2426 ( .A(n2833), .B(n2834), .C(n2835), .D(n2836), .S0(n3225), .S1(
        n3217), .Y(n2754) );
  MX4X1 U2427 ( .A(n2829), .B(n2830), .C(n2831), .D(n2832), .S0(n3225), .S1(
        n3217), .Y(n2755) );
  MX4X1 U2428 ( .A(n2821), .B(n2822), .C(n2823), .D(n2824), .S0(n3224), .S1(
        n3216), .Y(n2757) );
  NAND2X1 U2429 ( .A(n3771), .B(n465), .Y(MR) );
  CLKBUFX3 U2430 ( .A(n133), .Y(n3910) );
  CLKBUFX3 U2431 ( .A(n134), .Y(n3907) );
  CLKBUFX3 U2432 ( .A(n3185), .Y(n3188) );
  CLKBUFX3 U2433 ( .A(n3185), .Y(n3187) );
  NAND2X1 U2434 ( .A(n3659), .B(n3658), .Y(n3351) );
  NOR2X1 U2435 ( .A(n3657), .B(n3656), .Y(n3659) );
  MXI2X1 U2436 ( .A(n1522), .B(n3655), .S0(n3721), .Y(n3658) );
  NOR2X1 U2437 ( .A(n3749), .B(n3719), .Y(n3656) );
  NAND2X1 U2438 ( .A(n3664), .B(n3663), .Y(n3341) );
  NOR2X1 U2439 ( .A(n3662), .B(n3661), .Y(n3664) );
  MXI2X1 U2440 ( .A(n1523), .B(n3660), .S0(n3721), .Y(n3663) );
  NOR2X1 U2441 ( .A(n3749), .B(n3719), .Y(n3661) );
  NAND2X1 U2442 ( .A(n3131), .B(n3130), .Y(n2837) );
  NOR2X1 U2443 ( .A(n3129), .B(n3128), .Y(n3131) );
  MXI2X1 U2444 ( .A(n1524), .B(n3127), .S0(n3183), .Y(n3130) );
  NOR2X1 U2445 ( .A(n3212), .B(n3181), .Y(n3128) );
  NAND2X1 U2446 ( .A(n3669), .B(n3668), .Y(n3331) );
  NOR2X1 U2447 ( .A(n3667), .B(n3666), .Y(n3669) );
  MXI2X1 U2448 ( .A(n1524), .B(n3665), .S0(n3721), .Y(n3668) );
  NOR2X1 U2449 ( .A(n3749), .B(n3719), .Y(n3666) );
  NAND2X1 U2450 ( .A(n3136), .B(n3135), .Y(n2829) );
  NOR2X1 U2451 ( .A(n3134), .B(n3133), .Y(n3136) );
  MXI2X1 U2452 ( .A(n1525), .B(n3132), .S0(n3184), .Y(n3135) );
  NOR2X1 U2453 ( .A(n3212), .B(n3181), .Y(n3133) );
  NAND2X1 U2454 ( .A(n3674), .B(n3673), .Y(n3321) );
  NOR2X1 U2455 ( .A(n3672), .B(n3671), .Y(n3674) );
  MXI2X1 U2456 ( .A(n1525), .B(n3670), .S0(n3722), .Y(n3673) );
  NOR2X1 U2457 ( .A(n3749), .B(n3719), .Y(n3671) );
  NAND2X1 U2458 ( .A(n3141), .B(n3140), .Y(n2821) );
  NOR2X1 U2459 ( .A(n3139), .B(n3138), .Y(n3141) );
  MXI2X1 U2460 ( .A(n1526), .B(n3137), .S0(n3183), .Y(n3140) );
  NOR2X1 U2461 ( .A(n3212), .B(n3181), .Y(n3138) );
  NAND2X1 U2462 ( .A(n3679), .B(n3678), .Y(n3311) );
  NOR2X1 U2463 ( .A(n3677), .B(n3676), .Y(n3679) );
  MXI2X1 U2464 ( .A(n1526), .B(n3675), .S0(n3721), .Y(n3678) );
  NOR2X1 U2465 ( .A(n3749), .B(n3719), .Y(n3676) );
  NAND2X1 U2466 ( .A(n3684), .B(n3683), .Y(n3301) );
  NOR2X1 U2467 ( .A(n3682), .B(n3681), .Y(n3684) );
  MXI2X1 U2468 ( .A(n1527), .B(n3680), .S0(n3722), .Y(n3683) );
  NOR2X1 U2469 ( .A(n3749), .B(n3719), .Y(n3681) );
  CLKBUFX3 U2470 ( .A(n3185), .Y(n3186) );
  CLKINVX1 U2471 ( .A(n3214), .Y(n3190) );
  CLKINVX1 U2472 ( .A(n3214), .Y(n3189) );
  CLKBUFX3 U2473 ( .A(n3234), .Y(n3233) );
  CLKBUFX3 U2474 ( .A(n3234), .Y(n3232) );
  CLKBUFX3 U2475 ( .A(n136), .Y(n3899) );
  CLKBUFX3 U2476 ( .A(n137), .Y(n3896) );
  CLKBUFX3 U2477 ( .A(n138), .Y(n3893) );
  CLKBUFX3 U2478 ( .A(n139), .Y(n3890) );
  CLKBUFX3 U2479 ( .A(n140), .Y(n3887) );
  CLKBUFX3 U2480 ( .A(n141), .Y(n3884) );
  CLKBUFX3 U2481 ( .A(n136), .Y(n3900) );
  CLKBUFX3 U2482 ( .A(n137), .Y(n3897) );
  CLKBUFX3 U2483 ( .A(n138), .Y(n3894) );
  CLKBUFX3 U2484 ( .A(n139), .Y(n3891) );
  CLKBUFX3 U2485 ( .A(n140), .Y(n3888) );
  CLKBUFX3 U2486 ( .A(n141), .Y(n3885) );
  CLKBUFX3 U2487 ( .A(n3234), .Y(n3231) );
  CLKBUFX3 U2488 ( .A(n136), .Y(n3901) );
  CLKBUFX3 U2489 ( .A(n137), .Y(n3898) );
  CLKBUFX3 U2490 ( .A(n138), .Y(n3895) );
  CLKBUFX3 U2491 ( .A(n139), .Y(n3892) );
  CLKBUFX3 U2492 ( .A(n140), .Y(n3889) );
  CLKBUFX3 U2493 ( .A(n141), .Y(n3886) );
  CLKBUFX3 U2494 ( .A(n3222), .Y(n3220) );
  CLKBUFX3 U2495 ( .A(n3222), .Y(n3219) );
  CLKBUFX3 U2496 ( .A(n3222), .Y(n3218) );
  CLKBUFX3 U2497 ( .A(n3221), .Y(n3217) );
  CLKBUFX3 U2498 ( .A(n3221), .Y(n3216) );
  NAND2X1 U2499 ( .A(n3634), .B(n3633), .Y(n3401) );
  NOR2X1 U2500 ( .A(n3632), .B(n3631), .Y(n3634) );
  MXI2X1 U2501 ( .A(n1517), .B(n3630), .S0(n3720), .Y(n3633) );
  NOR2X1 U2502 ( .A(n3748), .B(n3719), .Y(n3631) );
  NAND2X1 U2503 ( .A(n3639), .B(n3638), .Y(n3391) );
  NOR2X1 U2504 ( .A(n3637), .B(n3636), .Y(n3639) );
  MXI2X1 U2505 ( .A(n1518), .B(n3635), .S0(n3720), .Y(n3638) );
  NOR2X1 U2506 ( .A(n3748), .B(n3719), .Y(n3636) );
  NAND2X1 U2507 ( .A(n3644), .B(n3643), .Y(n3381) );
  NOR2X1 U2508 ( .A(n3642), .B(n3641), .Y(n3644) );
  MXI2X1 U2509 ( .A(n1519), .B(n3640), .S0(n3721), .Y(n3643) );
  NOR2X1 U2510 ( .A(n3748), .B(n3719), .Y(n3641) );
  NAND2X1 U2511 ( .A(n3649), .B(n3648), .Y(n3371) );
  NOR2X1 U2512 ( .A(n3647), .B(n3646), .Y(n3649) );
  MXI2X1 U2513 ( .A(n1520), .B(n3645), .S0(n3721), .Y(n3648) );
  NOR2X1 U2514 ( .A(n3748), .B(n3719), .Y(n3646) );
  NAND2X1 U2515 ( .A(n3654), .B(n3653), .Y(n3361) );
  NOR2X1 U2516 ( .A(n3652), .B(n3651), .Y(n3654) );
  MXI2X1 U2517 ( .A(n1521), .B(n3650), .S0(n3721), .Y(n3653) );
  NOR2X1 U2518 ( .A(n3749), .B(n3719), .Y(n3651) );
  NAND2X1 U2519 ( .A(n3629), .B(n3628), .Y(n3411) );
  NOR2X1 U2520 ( .A(n3627), .B(n3626), .Y(n3629) );
  MXI2X1 U2521 ( .A(n1516), .B(n3625), .S0(n3721), .Y(n3628) );
  NOR2X1 U2522 ( .A(n3748), .B(n3719), .Y(n3626) );
  AND4X1 U2523 ( .A(n295), .B(n296), .C(n297), .D(n298), .Y(n121) );
  AOI221XL U2524 ( .A0(n299), .A1(n2693), .B0(N218), .B1(n300), .C0(n301), .Y(
        n298) );
  AOI222XL U2525 ( .A0(N788), .A1(n3782), .B0(N404), .B1(n250), .C0(N867), 
        .C1(n251), .Y(n296) );
  AOI222XL U2526 ( .A0(N436), .A1(n246), .B0(N660), .B1(n247), .C0(N596), .C1(
        n3780), .Y(n297) );
  CLKBUFX3 U2527 ( .A(n142), .Y(n3881) );
  CLKBUFX3 U2528 ( .A(n143), .Y(n3878) );
  CLKBUFX3 U2529 ( .A(n144), .Y(n3875) );
  CLKBUFX3 U2530 ( .A(n145), .Y(n3872) );
  CLKBUFX3 U2531 ( .A(n113), .Y(n3964) );
  CLKBUFX3 U2532 ( .A(n142), .Y(n3882) );
  CLKBUFX3 U2533 ( .A(n143), .Y(n3879) );
  CLKBUFX3 U2534 ( .A(n144), .Y(n3876) );
  CLKBUFX3 U2535 ( .A(n145), .Y(n3873) );
  CLKBUFX3 U2536 ( .A(n113), .Y(n3965) );
  AOI222XL U2537 ( .A0(N442), .A1(n246), .B0(N666), .B1(n247), .C0(N602), .C1(
        n248), .Y(n231) );
  CLKBUFX3 U2538 ( .A(n142), .Y(n3883) );
  CLKBUFX3 U2539 ( .A(n143), .Y(n3880) );
  CLKBUFX3 U2540 ( .A(n144), .Y(n3877) );
  CLKBUFX3 U2541 ( .A(n145), .Y(n3874) );
  CLKBUFX3 U2542 ( .A(n113), .Y(n3966) );
  NAND2X1 U2543 ( .A(n3604), .B(n3603), .Y(n3461) );
  NOR2X1 U2544 ( .A(n3602), .B(n3601), .Y(n3604) );
  MXI2X1 U2545 ( .A(n1511), .B(n3600), .S0(n3720), .Y(n3603) );
  NOR2X1 U2546 ( .A(n3747), .B(n3720), .Y(n3601) );
  NAND2X1 U2547 ( .A(n3609), .B(n3608), .Y(n3451) );
  NOR2X1 U2548 ( .A(n3607), .B(n3606), .Y(n3609) );
  MXI2X1 U2549 ( .A(n1512), .B(n3605), .S0(n3720), .Y(n3608) );
  NOR2X1 U2550 ( .A(n3747), .B(n3719), .Y(n3606) );
  NAND2X1 U2551 ( .A(n3614), .B(n3613), .Y(n3441) );
  NOR2X1 U2552 ( .A(n3612), .B(n3611), .Y(n3614) );
  MXI2X1 U2553 ( .A(n1513), .B(n3610), .S0(n3720), .Y(n3613) );
  NOR2X1 U2554 ( .A(n3747), .B(n3719), .Y(n3611) );
  NAND2X1 U2555 ( .A(n3619), .B(n3618), .Y(n3431) );
  NOR2X1 U2556 ( .A(n3617), .B(n3616), .Y(n3619) );
  MXI2X1 U2557 ( .A(n1514), .B(n3615), .S0(n3720), .Y(n3618) );
  NOR2X1 U2558 ( .A(n3747), .B(n3719), .Y(n3616) );
  NAND2X1 U2559 ( .A(n3624), .B(n3623), .Y(n3421) );
  NOR2X1 U2560 ( .A(n3622), .B(n3621), .Y(n3624) );
  MXI2X1 U2561 ( .A(n1515), .B(n3620), .S0(n3720), .Y(n3623) );
  NOR2X1 U2562 ( .A(n3748), .B(n3719), .Y(n3621) );
  AND2X2 U2563 ( .A(N87), .B(n3973), .Y(N153) );
  AND2X2 U2564 ( .A(N90), .B(n3973), .Y(N156) );
  AND2X2 U2565 ( .A(N85), .B(n3973), .Y(N151) );
  AND2X2 U2566 ( .A(N86), .B(n3973), .Y(N152) );
  AND2X2 U2567 ( .A(N89), .B(n3973), .Y(N155) );
  AND2X2 U2568 ( .A(N84), .B(n3973), .Y(N150) );
  AND2X2 U2569 ( .A(N88), .B(n3973), .Y(N154) );
  AOI221XL U2570 ( .A0(N960), .A1(n470), .B0(n471), .B1(n4024), .C0(n472), .Y(
        n469) );
  OAI221XL U2571 ( .A0(n3787), .A1(n244), .B0(n4039), .B1(n3792), .C0(n245), 
        .Y(n471) );
  OAI2BB2XL U2572 ( .B0(n3787), .B1(n237), .A0N(n473), .A1N(n2670), .Y(n472)
         );
  AND4X1 U2573 ( .A(n287), .B(n288), .C(n289), .D(n290), .Y(n120) );
  AOI221XL U2574 ( .A0(n291), .A1(n2686), .B0(N217), .B1(n292), .C0(n293), .Y(
        n290) );
  AOI222XL U2575 ( .A0(N789), .A1(n249), .B0(N405), .B1(n250), .C0(N868), .C1(
        n251), .Y(n288) );
  AOI222XL U2576 ( .A0(N437), .A1(n3774), .B0(N661), .B1(n3781), .C0(N597), 
        .C1(n248), .Y(n289) );
  AND4X1 U2577 ( .A(n317), .B(n318), .C(n319), .D(n320), .Y(n124) );
  AOI221XL U2578 ( .A0(n321), .A1(n2683), .B0(N219), .B1(n322), .C0(n323), .Y(
        n320) );
  AOI222XL U2579 ( .A0(N787), .A1(n249), .B0(N403), .B1(n250), .C0(N866), .C1(
        n251), .Y(n318) );
  AOI222XL U2580 ( .A0(N435), .A1(n3774), .B0(N659), .B1(n3781), .C0(N595), 
        .C1(n248), .Y(n319) );
  AND4X1 U2581 ( .A(n385), .B(n386), .C(n387), .D(n388), .Y(n135) );
  AOI222XL U2582 ( .A0(N786), .A1(n3782), .B0(N402), .B1(n250), .C0(N865), 
        .C1(n251), .Y(n386) );
  AOI222XL U2583 ( .A0(N434), .A1(n246), .B0(N658), .B1(n247), .C0(N594), .C1(
        n3780), .Y(n387) );
  AOI221XL U2584 ( .A0(n389), .A1(n4023), .B0(N220), .B1(n390), .C0(n391), .Y(
        n388) );
  CLKBUFX3 U2585 ( .A(n116), .Y(n3959) );
  CLKBUFX3 U2586 ( .A(n117), .Y(n3956) );
  CLKBUFX3 U2587 ( .A(n118), .Y(n3953) );
  CLKBUFX3 U2588 ( .A(n119), .Y(n3950) );
  CLKBUFX3 U2589 ( .A(n146), .Y(n3870) );
  CLKBUFX3 U2590 ( .A(n116), .Y(n3960) );
  CLKBUFX3 U2591 ( .A(n117), .Y(n3957) );
  CLKBUFX3 U2592 ( .A(n118), .Y(n3954) );
  CLKBUFX3 U2593 ( .A(n119), .Y(n3951) );
  CLKBUFX3 U2594 ( .A(n146), .Y(n3869) );
  CLKINVX1 U2595 ( .A(n513), .Y(n3993) );
  OAI31XL U2596 ( .A0(n514), .A1(n515), .A2(n516), .B0(n4045), .Y(n513) );
  OA22X1 U2597 ( .A0(n4008), .A1(n518), .B0(n519), .B1(n520), .Y(n514) );
  AOI222XL U2598 ( .A0(N441), .A1(n3774), .B0(N665), .B1(n247), .C0(N601), 
        .C1(n248), .Y(n257) );
  AOI222XL U2599 ( .A0(N440), .A1(n246), .B0(N664), .B1(n247), .C0(N600), .C1(
        n248), .Y(n265) );
  AOI222XL U2600 ( .A0(N439), .A1(n3774), .B0(N663), .B1(n247), .C0(N599), 
        .C1(n248), .Y(n273) );
  AOI222XL U2601 ( .A0(N438), .A1(n246), .B0(N662), .B1(n247), .C0(N598), .C1(
        n248), .Y(n281) );
  CLKBUFX3 U2602 ( .A(n146), .Y(n3871) );
  CLKBUFX3 U2603 ( .A(n116), .Y(n3961) );
  CLKBUFX3 U2604 ( .A(n117), .Y(n3958) );
  CLKBUFX3 U2605 ( .A(n118), .Y(n3955) );
  CLKBUFX3 U2606 ( .A(n119), .Y(n3952) );
  NAND2X1 U2607 ( .A(n3594), .B(n3593), .Y(n3481) );
  NOR2X1 U2608 ( .A(n3592), .B(n3591), .Y(n3594) );
  MXI2X1 U2609 ( .A(n1509), .B(n3590), .S0(n3720), .Y(n3593) );
  NOR2X1 U2610 ( .A(n3747), .B(n3720), .Y(n3591) );
  NAND2X1 U2611 ( .A(n3559), .B(n3558), .Y(n3551) );
  NOR2X1 U2612 ( .A(n3557), .B(n3556), .Y(n3559) );
  MXI2X1 U2613 ( .A(n1502), .B(n3555), .S0(n3722), .Y(n3558) );
  NOR2X1 U2614 ( .A(n3746), .B(n3720), .Y(n3556) );
  NAND2X1 U2615 ( .A(n3564), .B(n3563), .Y(n3541) );
  NOR2X1 U2616 ( .A(n3562), .B(n3561), .Y(n3564) );
  MXI2X1 U2617 ( .A(n1503), .B(n3560), .S0(n3722), .Y(n3563) );
  NOR2X1 U2618 ( .A(n3746), .B(n3720), .Y(n3561) );
  NAND2X1 U2619 ( .A(n3569), .B(n3568), .Y(n3531) );
  NOR2X1 U2620 ( .A(n3567), .B(n3566), .Y(n3569) );
  MXI2X1 U2621 ( .A(n1504), .B(n3565), .S0(n3722), .Y(n3568) );
  NOR2X1 U2622 ( .A(n3746), .B(n3720), .Y(n3566) );
  NAND2X1 U2623 ( .A(n3574), .B(n3573), .Y(n3521) );
  NOR2X1 U2624 ( .A(n3572), .B(n3571), .Y(n3574) );
  MXI2X1 U2625 ( .A(n1505), .B(n3570), .S0(n3722), .Y(n3573) );
  NOR2X1 U2626 ( .A(n3746), .B(n3720), .Y(n3571) );
  NAND2X1 U2627 ( .A(n3579), .B(n3578), .Y(n3511) );
  NOR2X1 U2628 ( .A(n3577), .B(n3576), .Y(n3579) );
  MXI2X1 U2629 ( .A(n1506), .B(n3575), .S0(n3721), .Y(n3578) );
  NOR2X1 U2630 ( .A(n3746), .B(n3720), .Y(n3576) );
  NAND2X1 U2631 ( .A(n3584), .B(n3583), .Y(n3501) );
  NOR2X1 U2632 ( .A(n3582), .B(n3581), .Y(n3584) );
  MXI2X1 U2633 ( .A(n1507), .B(n3580), .S0(n3721), .Y(n3583) );
  NOR2X1 U2634 ( .A(n3746), .B(n3720), .Y(n3581) );
  NAND2X1 U2635 ( .A(n3589), .B(n3588), .Y(n3491) );
  NOR2X1 U2636 ( .A(n3587), .B(n3586), .Y(n3589) );
  MXI2X1 U2637 ( .A(n1508), .B(n3585), .S0(n3721), .Y(n3588) );
  NOR2X1 U2638 ( .A(n3747), .B(n3720), .Y(n3586) );
  NAND2X1 U2639 ( .A(n3599), .B(n3598), .Y(n3471) );
  NOR2X1 U2640 ( .A(n3597), .B(n3596), .Y(n3599) );
  MXI2X1 U2641 ( .A(n1510), .B(n3595), .S0(n3721), .Y(n3598) );
  NOR2X1 U2642 ( .A(n3747), .B(n3720), .Y(n3596) );
  AND2X2 U2643 ( .A(N79), .B(n3973), .Y(N145) );
  AND2X2 U2644 ( .A(N83), .B(n3973), .Y(N149) );
  AND2X2 U2645 ( .A(N77), .B(n3973), .Y(N143) );
  AND2X2 U2646 ( .A(N78), .B(n3973), .Y(N144) );
  AND2X2 U2647 ( .A(N81), .B(n3973), .Y(N147) );
  AND2X2 U2648 ( .A(N82), .B(n3973), .Y(N148) );
  AND2X2 U2649 ( .A(N80), .B(n3973), .Y(N146) );
  OAI22XL U2650 ( .A0(n3996), .A1(n4025), .B0(n3972), .B1(n237), .Y(n429) );
  OAI22XL U2651 ( .A0(n3996), .A1(n4026), .B0(n3978), .B1(n237), .Y(n437) );
  OAI22XL U2652 ( .A0(n3996), .A1(n4027), .B0(n3979), .B1(n237), .Y(n445) );
  OAI22XL U2653 ( .A0(n3996), .A1(n4028), .B0(n3981), .B1(n237), .Y(n453) );
  OAI22XL U2654 ( .A0(n3996), .A1(n4029), .B0(n3982), .B1(n237), .Y(n461) );
  OAI22XL U2655 ( .A0(n3996), .A1(n4030), .B0(n4040), .B1(n237), .Y(n235) );
  OAI22XL U2656 ( .A0(n3996), .A1(n4031), .B0(n4041), .B1(n237), .Y(n261) );
  OAI22XL U2657 ( .A0(n3996), .A1(n4032), .B0(n4042), .B1(n237), .Y(n269) );
  OAI22XL U2658 ( .A0(n3996), .A1(n4033), .B0(n4043), .B1(n237), .Y(n277) );
  OAI22XL U2659 ( .A0(n3996), .A1(n4034), .B0(n4044), .B1(n237), .Y(n285) );
  OAI22XL U2660 ( .A0(n3996), .A1(n4035), .B0(n3977), .B1(n237), .Y(n293) );
  OAI22XL U2661 ( .A0(n3996), .A1(n4036), .B0(n3976), .B1(n237), .Y(n301) );
  OAI22XL U2662 ( .A0(n3996), .A1(n4037), .B0(n3975), .B1(n237), .Y(n323) );
  OAI22XL U2663 ( .A0(n3996), .A1(n4038), .B0(n3974), .B1(n237), .Y(n391) );
  NAND2X1 U2664 ( .A(n158), .B(n148), .Y(n228) );
  AND2X2 U2665 ( .A(n180), .B(n164), .Y(n216) );
  AND2X2 U2666 ( .A(n179), .B(n180), .Y(n170) );
  AND2X2 U2667 ( .A(n179), .B(n190), .Y(n183) );
  AND2X2 U2668 ( .A(n179), .B(n163), .Y(n193) );
  AND2X2 U2669 ( .A(n179), .B(n203), .Y(n206) );
  AND2X2 U2670 ( .A(n163), .B(n164), .Y(n155) );
  AND2X2 U2671 ( .A(n164), .B(n190), .Y(n148) );
  NAND2X1 U2672 ( .A(n147), .B(n148), .Y(n114) );
  NOR3X1 U2673 ( .A(n464), .B(n3973), .C(n465), .Y(n213) );
  NAND2X1 U2674 ( .A(n151), .B(n148), .Y(n149) );
  AND2X2 U2675 ( .A(n521), .B(n4045), .Y(n480) );
  NAND4X1 U2676 ( .A(n464), .B(n3995), .C(n523), .D(n111), .Y(n521) );
  OAI22XL U2677 ( .A0(n519), .A1(n4008), .B0(n518), .B1(n520), .Y(n523) );
  AND2X2 U2678 ( .A(n203), .B(n164), .Y(n167) );
  NAND2X1 U2679 ( .A(n170), .B(n147), .Y(n175) );
  NAND2X1 U2680 ( .A(n183), .B(n147), .Y(n186) );
  NAND2X1 U2681 ( .A(n193), .B(n147), .Y(n196) );
  NAND2X1 U2682 ( .A(n206), .B(n147), .Y(n209) );
  NAND2X1 U2683 ( .A(n216), .B(n147), .Y(n219) );
  NAND2X1 U2684 ( .A(n155), .B(n147), .Y(n159) );
  NAND2X1 U2685 ( .A(n167), .B(n147), .Y(n201) );
  OAI21XL U2686 ( .A0(N226), .A1(n3792), .B0(n2656), .Y(n341) );
  OAI21XL U2687 ( .A0(N228), .A1(n3792), .B0(n2656), .Y(n353) );
  OAI21XL U2688 ( .A0(N230), .A1(n3792), .B0(n2656), .Y(n365) );
  OAI21XL U2689 ( .A0(N232), .A1(n3791), .B0(n2656), .Y(n377) );
  OAI21XL U2690 ( .A0(N234), .A1(n3791), .B0(n2656), .Y(n397) );
  OAI21XL U2691 ( .A0(N238), .A1(n3791), .B0(n2656), .Y(n421) );
  OAI21XL U2692 ( .A0(N223), .A1(n3791), .B0(n2656), .Y(n315) );
  OAI21XL U2693 ( .A0(N227), .A1(n3792), .B0(n2656), .Y(n347) );
  OAI21XL U2694 ( .A0(N229), .A1(n3791), .B0(n2656), .Y(n359) );
  OAI21XL U2695 ( .A0(N231), .A1(n3792), .B0(n2656), .Y(n371) );
  OAI21XL U2696 ( .A0(N233), .A1(n3791), .B0(n2656), .Y(n383) );
  OAI21XL U2697 ( .A0(N235), .A1(n3791), .B0(n2656), .Y(n403) );
  OAI21XL U2698 ( .A0(N236), .A1(n3791), .B0(n2656), .Y(n409) );
  OAI21XL U2699 ( .A0(N237), .A1(n3791), .B0(n2656), .Y(n415) );
  NAND2X1 U2700 ( .A(n170), .B(n151), .Y(n177) );
  NAND2X1 U2701 ( .A(n183), .B(n151), .Y(n188) );
  NAND2X1 U2702 ( .A(n193), .B(n151), .Y(n198) );
  NAND2X1 U2703 ( .A(n206), .B(n151), .Y(n211) );
  NAND2X1 U2704 ( .A(n216), .B(n151), .Y(n222) );
  NAND2X1 U2705 ( .A(n155), .B(n151), .Y(n161) );
  OAI21XL U2706 ( .A0(N225), .A1(n3791), .B0(n2656), .Y(n335) );
  OAI21XL U2707 ( .A0(N224), .A1(n3791), .B0(n2656), .Y(n329) );
  OAI21XL U2708 ( .A0(N222), .A1(n3791), .B0(n2656), .Y(n307) );
  NAND2X1 U2709 ( .A(n170), .B(n154), .Y(n168) );
  NAND2X1 U2710 ( .A(n170), .B(n158), .Y(n171) );
  NAND2X1 U2711 ( .A(n183), .B(n154), .Y(n181) );
  NAND2X1 U2712 ( .A(n183), .B(n158), .Y(n184) );
  NAND2X1 U2713 ( .A(n193), .B(n154), .Y(n191) );
  NAND2X1 U2714 ( .A(n193), .B(n158), .Y(n194) );
  NAND2X1 U2715 ( .A(n206), .B(n154), .Y(n204) );
  NAND2X1 U2716 ( .A(n206), .B(n158), .Y(n207) );
  NAND2X1 U2717 ( .A(n216), .B(n154), .Y(n214) );
  NAND2X1 U2718 ( .A(n216), .B(n158), .Y(n217) );
  NAND2X1 U2719 ( .A(n167), .B(n154), .Y(n165) );
  NAND2X1 U2720 ( .A(n167), .B(n158), .Y(n173) );
  NAND2X1 U2721 ( .A(n154), .B(n148), .Y(n225) );
  NAND2X1 U2722 ( .A(n154), .B(n155), .Y(n152) );
  NAND2X1 U2723 ( .A(n158), .B(n155), .Y(n156) );
  CLKINVX1 U2724 ( .A(N239), .Y(n4025) );
  CLKINVX1 U2725 ( .A(N240), .Y(n4026) );
  CLKINVX1 U2726 ( .A(N248), .Y(n4034) );
  OAI221XL U2727 ( .A0(n238), .A1(n4039), .B0(n3792), .B1(N253), .C0(n474), 
        .Y(n473) );
  AOI221XL U2728 ( .A0(N656), .A1(n242), .B0(n3787), .B1(n3998), .C0(n243), 
        .Y(n474) );
  AO22X1 U2729 ( .A0(N401), .A1(n250), .B0(N433), .B1(n246), .Y(n477) );
  OAI221XL U2730 ( .A0(n3978), .A1(n244), .B0(n4026), .B1(n3793), .C0(n245), 
        .Y(n435) );
  OAI221XL U2731 ( .A0(n3979), .A1(n244), .B0(n4027), .B1(n3793), .C0(n245), 
        .Y(n443) );
  OAI221XL U2732 ( .A0(n3981), .A1(n244), .B0(n4028), .B1(n3793), .C0(n245), 
        .Y(n451) );
  OAI221XL U2733 ( .A0(n3982), .A1(n244), .B0(n4029), .B1(n3793), .C0(n245), 
        .Y(n459) );
  OAI221XL U2734 ( .A0(n4040), .A1(n244), .B0(n4030), .B1(n3792), .C0(n245), 
        .Y(n233) );
  OAI221XL U2735 ( .A0(n4041), .A1(n244), .B0(n4031), .B1(n3792), .C0(n245), 
        .Y(n259) );
  OAI221XL U2736 ( .A0(n4044), .A1(n244), .B0(n4034), .B1(n3792), .C0(n245), 
        .Y(n283) );
  OAI221XL U2737 ( .A0(n3977), .A1(n244), .B0(n4035), .B1(n3792), .C0(n245), 
        .Y(n291) );
  OAI221XL U2738 ( .A0(n3974), .A1(n244), .B0(n4038), .B1(n3792), .C0(n245), 
        .Y(n389) );
  OAI221XL U2739 ( .A0(n3972), .A1(n244), .B0(n4025), .B1(n3792), .C0(n245), 
        .Y(n427) );
  OAI221XL U2740 ( .A0(n4043), .A1(n244), .B0(n4033), .B1(n3792), .C0(n245), 
        .Y(n275) );
  OAI221XL U2741 ( .A0(n3976), .A1(n244), .B0(n4036), .B1(n3792), .C0(n245), 
        .Y(n299) );
  OAI221XL U2742 ( .A0(n3975), .A1(n244), .B0(n4037), .B1(n3792), .C0(n245), 
        .Y(n321) );
  OAI221XL U2743 ( .A0(n4042), .A1(n244), .B0(n4032), .B1(n3792), .C0(n245), 
        .Y(n267) );
  OAI221XL U2744 ( .A0(n4038), .A1(n238), .B0(N252), .B1(n3792), .C0(n392), 
        .Y(n390) );
  AOI221XL U2745 ( .A0(n3998), .A1(n3974), .B0(n242), .B1(instruction[1]), 
        .C0(n243), .Y(n392) );
  OAI221XL U2746 ( .A0(n4026), .A1(n3773), .B0(N240), .B1(n3792), .C0(n438), 
        .Y(n436) );
  AOI221XL U2747 ( .A0(n3998), .A1(n3978), .B0(n242), .B1(N54), .C0(n243), .Y(
        n438) );
  OAI221XL U2748 ( .A0(n4028), .A1(n3773), .B0(N242), .B1(n3793), .C0(n454), 
        .Y(n452) );
  AOI221XL U2749 ( .A0(n3998), .A1(n3981), .B0(n242), .B1(n3980), .C0(n243), 
        .Y(n454) );
  OAI221XL U2750 ( .A0(n4029), .A1(n238), .B0(N243), .B1(n3793), .C0(n463), 
        .Y(n460) );
  AOI221XL U2751 ( .A0(n3998), .A1(n3982), .B0(n242), .B1(N51), .C0(n243), .Y(
        n463) );
  OAI221XL U2752 ( .A0(n4035), .A1(n3773), .B0(N249), .B1(n3792), .C0(n294), 
        .Y(n292) );
  AOI221XL U2753 ( .A0(n3998), .A1(n3977), .B0(n242), .B1(instruction[4]), 
        .C0(n243), .Y(n294) );
  OAI221XL U2754 ( .A0(n4027), .A1(n238), .B0(N241), .B1(n3793), .C0(n446), 
        .Y(n444) );
  AOI221XL U2755 ( .A0(n3998), .A1(n3979), .B0(n242), .B1(N53), .C0(n243), .Y(
        n446) );
  OAI221XL U2756 ( .A0(n4025), .A1(n238), .B0(N239), .B1(n3792), .C0(n430), 
        .Y(n428) );
  AOI221XL U2757 ( .A0(n3998), .A1(n3972), .B0(n242), .B1(\seIM[31] ), .C0(
        n243), .Y(n430) );
  OAI221XL U2758 ( .A0(n4036), .A1(n238), .B0(N250), .B1(n3792), .C0(n302), 
        .Y(n300) );
  AOI221XL U2759 ( .A0(n3998), .A1(n3976), .B0(n242), .B1(instruction[3]), 
        .C0(n243), .Y(n302) );
  OAI221XL U2760 ( .A0(n4037), .A1(n3773), .B0(N251), .B1(n3792), .C0(n324), 
        .Y(n322) );
  AOI221XL U2761 ( .A0(n3998), .A1(n3975), .B0(n242), .B1(instruction[2]), 
        .C0(n243), .Y(n324) );
  AND2X2 U2762 ( .A(N69), .B(n3973), .Y(N135) );
  AND2X2 U2763 ( .A(N75), .B(n3973), .Y(N141) );
  AND2X2 U2764 ( .A(N71), .B(n3973), .Y(N137) );
  AND2X2 U2765 ( .A(N73), .B(n3973), .Y(N139) );
  AND2X2 U2766 ( .A(N74), .B(n3973), .Y(N140) );
  AND2X2 U2767 ( .A(N72), .B(n3973), .Y(N138) );
  AND2X2 U2768 ( .A(N76), .B(n3973), .Y(N142) );
  AND2X2 U2769 ( .A(N70), .B(n3973), .Y(N136) );
  NAND2X1 U2770 ( .A(n536), .B(n4045), .Y(n3783) );
  NAND2X1 U2771 ( .A(n536), .B(n4045), .Y(n478) );
  AND2X2 U2772 ( .A(N61), .B(n3973), .Y(N127) );
  AND2X2 U2773 ( .A(N65), .B(n3973), .Y(N131) );
  AND2X2 U2774 ( .A(N62), .B(n3973), .Y(N128) );
  AND2X2 U2775 ( .A(N63), .B(n3973), .Y(N129) );
  AND2X2 U2776 ( .A(N64), .B(n3973), .Y(N130) );
  AND2X2 U2777 ( .A(N67), .B(n3973), .Y(N133) );
  AND2X2 U2778 ( .A(N68), .B(n3973), .Y(N134) );
  AND2X2 U2779 ( .A(N66), .B(n3973), .Y(N132) );
  AND2X2 U2780 ( .A(n563), .B(n3999), .Y(n554) );
  NAND3X1 U2781 ( .A(n237), .B(n475), .C(n559), .Y(n243) );
  NAND3X1 U2782 ( .A(n552), .B(n3999), .C(n540), .Y(n559) );
  AND4X1 U2783 ( .A(n547), .B(n548), .C(n549), .D(n550), .Y(n464) );
  NOR4X1 U2784 ( .A(n254), .B(n3777), .C(n3778), .D(n3779), .Y(n548) );
  NOR4BX1 U2785 ( .AN(n2656), .B(n3780), .C(n3781), .D(n252), .Y(n549) );
  NOR4BX1 U2786 ( .AN(n476), .B(n3997), .C(n470), .D(n3782), .Y(n550) );
  NAND2X1 U2787 ( .A(n551), .B(n554), .Y(n239) );
  NAND2X1 U2788 ( .A(n561), .B(n551), .Y(n244) );
  NAND2X1 U2789 ( .A(n560), .B(n554), .Y(n475) );
  NAND2X1 U2790 ( .A(n475), .B(n476), .Y(n462) );
  AND2X2 U2791 ( .A(n562), .B(n551), .Y(n250) );
  NAND2X1 U2792 ( .A(n554), .B(n525), .Y(n3773) );
  NAND2X1 U2793 ( .A(n554), .B(n525), .Y(n238) );
  AND2X2 U2794 ( .A(n562), .B(n551), .Y(n3779) );
  AND2X2 U2795 ( .A(n553), .B(n554), .Y(n3777) );
  AND2X2 U2796 ( .A(n553), .B(n554), .Y(n253) );
  NAND4X1 U2797 ( .A(n464), .B(n3995), .C(n537), .D(n538), .Y(MW) );
  NOR2X1 U2798 ( .A(n516), .B(n465), .Y(n537) );
  NOR4X1 U2799 ( .A(n536), .B(n519), .C(n518), .D(n515), .Y(n538) );
  AND2X2 U2800 ( .A(n561), .B(n525), .Y(n242) );
  AND2X2 U2801 ( .A(n553), .B(n524), .Y(n247) );
  AND2X2 U2802 ( .A(n553), .B(n524), .Y(n3781) );
  AND2X2 U2803 ( .A(n562), .B(n553), .Y(n3774) );
  AND2X2 U2804 ( .A(n551), .B(n524), .Y(n248) );
  AND2X2 U2805 ( .A(n540), .B(n543), .Y(n519) );
  CLKINVX1 U2806 ( .A(n245), .Y(n3997) );
  AND2X2 U2807 ( .A(n539), .B(n3999), .Y(n252) );
  AND3X2 U2808 ( .A(n552), .B(n3999), .C(n3994), .Y(n562) );
  NOR2X1 U2809 ( .A(n4006), .B(n4005), .Y(n180) );
  AND2X2 U2810 ( .A(n539), .B(n3999), .Y(n3772) );
  NOR2BX1 U2811 ( .AN(N238), .B(n3971), .Y(datain[15]) );
  NOR2BX1 U2812 ( .AN(N237), .B(n3971), .Y(datain[16]) );
  NOR2BX1 U2813 ( .AN(N236), .B(n3971), .Y(datain[17]) );
  NOR2BX1 U2814 ( .AN(N235), .B(n3971), .Y(datain[18]) );
  NOR2BX1 U2815 ( .AN(N234), .B(n3971), .Y(datain[19]) );
  NOR2BX1 U2816 ( .AN(N233), .B(n3971), .Y(datain[20]) );
  NOR2BX1 U2817 ( .AN(N232), .B(n3971), .Y(datain[21]) );
  NOR2BX1 U2818 ( .AN(N231), .B(n3971), .Y(datain[22]) );
  NOR2BX1 U2819 ( .AN(N230), .B(n3971), .Y(datain[23]) );
  NOR2BX1 U2820 ( .AN(N229), .B(n3971), .Y(datain[24]) );
  NOR2BX1 U2821 ( .AN(N228), .B(n3971), .Y(datain[25]) );
  NOR2BX1 U2822 ( .AN(N227), .B(n3971), .Y(datain[26]) );
  NOR2BX1 U2823 ( .AN(N226), .B(n3971), .Y(datain[27]) );
  NOR2BX1 U2824 ( .AN(N225), .B(n3971), .Y(datain[28]) );
  NOR2BX1 U2825 ( .AN(N224), .B(n3971), .Y(datain[29]) );
  NOR2BX1 U2826 ( .AN(N223), .B(n3971), .Y(datain[30]) );
  NOR2BX1 U2827 ( .AN(N222), .B(n3971), .Y(datain[31]) );
  OAI22XL U2828 ( .A0(n3941), .A1(n3851), .B0(n574), .B1(n3852), .Y(n1608) );
  OAI22XL U2829 ( .A0(n3941), .A1(n3849), .B0(n606), .B1(n3850), .Y(n1640) );
  OAI22XL U2830 ( .A0(n3941), .A1(n3844), .B0(n638), .B1(n3845), .Y(n1672) );
  OAI22XL U2831 ( .A0(n3941), .A1(n3842), .B0(n670), .B1(n3843), .Y(n1704) );
  OAI22XL U2832 ( .A0(n3942), .A1(n3839), .B0(n702), .B1(n3840), .Y(n1736) );
  OAI22XL U2833 ( .A0(n3942), .A1(n3837), .B0(n734), .B1(n3838), .Y(n1768) );
  OAI22XL U2834 ( .A0(n3942), .A1(n3835), .B0(n766), .B1(n3836), .Y(n1800) );
  OAI22XL U2835 ( .A0(n3942), .A1(n3833), .B0(n798), .B1(n3834), .Y(n1832) );
  OAI22XL U2836 ( .A0(n3942), .A1(n3830), .B0(n830), .B1(n3831), .Y(n1864) );
  OAI22XL U2837 ( .A0(n3942), .A1(n3828), .B0(n862), .B1(n3829), .Y(n1896) );
  OAI22XL U2838 ( .A0(n3942), .A1(n3826), .B0(n894), .B1(n3827), .Y(n1928) );
  OAI22XL U2839 ( .A0(n3942), .A1(n3824), .B0(n926), .B1(n3825), .Y(n1960) );
  OAI22XL U2840 ( .A0(n3942), .A1(n3819), .B0(n958), .B1(n3820), .Y(n1992) );
  OAI22XL U2841 ( .A0(n3942), .A1(n3817), .B0(n990), .B1(n3818), .Y(n2024) );
  OAI22XL U2842 ( .A0(n3942), .A1(n3815), .B0(n1022), .B1(n3816), .Y(n2056) );
  OAI22XL U2843 ( .A0(n3943), .A1(n3813), .B0(n1054), .B1(n3814), .Y(n2088) );
  OAI22XL U2844 ( .A0(n3943), .A1(n3809), .B0(n1086), .B1(n3810), .Y(n2120) );
  OAI22XL U2845 ( .A0(n3943), .A1(n3806), .B0(n1118), .B1(n3807), .Y(n2152) );
  OAI22XL U2846 ( .A0(n3943), .A1(n3804), .B0(n1150), .B1(n3805), .Y(n2184) );
  OAI22XL U2847 ( .A0(n3943), .A1(n3801), .B0(n1182), .B1(n3802), .Y(n2216) );
  OAI22XL U2848 ( .A0(n3943), .A1(n3799), .B0(n1214), .B1(n3800), .Y(n2248) );
  OAI22XL U2849 ( .A0(n3941), .A1(n3962), .B0(n1278), .B1(n3963), .Y(n2312) );
  OAI22XL U2850 ( .A0(n3941), .A1(n3867), .B0(n1310), .B1(n3868), .Y(n2344) );
  OAI22XL U2851 ( .A0(n3941), .A1(n3864), .B0(n1342), .B1(n3865), .Y(n2376) );
  OAI22XL U2852 ( .A0(n3941), .A1(n3861), .B0(n1374), .B1(n3862), .Y(n2408) );
  OAI22XL U2853 ( .A0(n3941), .A1(n3858), .B0(n1406), .B1(n3859), .Y(n2440) );
  OAI22XL U2854 ( .A0(n3941), .A1(n3855), .B0(n1438), .B1(n3856), .Y(n2472) );
  OAI22XL U2855 ( .A0(n3941), .A1(n3853), .B0(n1470), .B1(n3854), .Y(n2504) );
  OAI22XL U2856 ( .A0(n3941), .A1(n3847), .B0(n1502), .B1(n3848), .Y(n2536) );
  OAI22XL U2857 ( .A0(n3942), .A1(n3821), .B0(n1534), .B1(n3822), .Y(n2568) );
  AOI222XL U2858 ( .A0(dataout[31]), .A1(n3772), .B0(N959), .B1(n3775), .C0(
        n3997), .C1(n2735), .Y(n303) );
  NOR2X1 U2859 ( .A(\R[3][1] ), .B(n3204), .Y(n3167) );
  MXI4X1 U2860 ( .A(\R[20][1] ), .B(\R[21][1] ), .C(\R[22][1] ), .D(\R[23][1] ), .S0(n3179), .S1(n3206), .Y(n2771) );
  MXI4X1 U2861 ( .A(\R[4][1] ), .B(\R[5][1] ), .C(\R[6][1] ), .D(\R[7][1] ), 
        .S0(n3179), .S1(n3206), .Y(n2775) );
  MXI4X1 U2862 ( .A(\R[16][1] ), .B(\R[17][1] ), .C(\R[18][1] ), .D(\R[19][1] ), .S0(n3179), .S1(n3206), .Y(n2769) );
  MXI4X1 U2863 ( .A(\R[24][1] ), .B(\R[25][1] ), .C(\R[26][1] ), .D(\R[27][1] ), .S0(n3179), .S1(n3206), .Y(n2770) );
  MXI4X1 U2864 ( .A(\R[8][1] ), .B(\R[9][1] ), .C(\R[10][1] ), .D(\R[11][1] ), 
        .S0(n3179), .S1(n3206), .Y(n2774) );
  MXI4X1 U2865 ( .A(\R[28][1] ), .B(\R[29][1] ), .C(\R[30][1] ), .D(\R[31][1] ), .S0(n3179), .S1(n3206), .Y(n2772) );
  CLKMX2X2 U2866 ( .A(n3280), .B(n3275), .S0(n3767), .Y(N249) );
  MXI4X1 U2867 ( .A(n3281), .B(n3282), .C(n3283), .D(n3284), .S0(n3760), .S1(
        n3752), .Y(n3280) );
  MXI4X1 U2868 ( .A(n3276), .B(n3277), .C(n3278), .D(n3279), .S0(n3760), .S1(
        n3752), .Y(n3275) );
  MXI4X1 U2869 ( .A(\R[12][4] ), .B(\R[13][4] ), .C(\R[14][4] ), .D(\R[15][4] ), .S0(n3717), .S1(n3743), .Y(n3284) );
  MXI4X1 U2870 ( .A(n3286), .B(n3287), .C(n3288), .D(n3289), .S0(n3760), .S1(
        n3752), .Y(n3285) );
  OAI22XL U2871 ( .A0(n3938), .A1(n3851), .B0(n575), .B1(n3852), .Y(n1609) );
  OAI22XL U2872 ( .A0(n3932), .A1(n3851), .B0(n576), .B1(n3852), .Y(n1610) );
  OAI22XL U2873 ( .A0(n3929), .A1(n168), .B0(n577), .B1(n3852), .Y(n1611) );
  OAI22XL U2874 ( .A0(n3926), .A1(n168), .B0(n578), .B1(n3852), .Y(n1612) );
  OAI22XL U2875 ( .A0(n3923), .A1(n3851), .B0(n579), .B1(n3852), .Y(n1613) );
  OAI22XL U2876 ( .A0(n3938), .A1(n3849), .B0(n607), .B1(n3850), .Y(n1641) );
  OAI22XL U2877 ( .A0(n3932), .A1(n3849), .B0(n608), .B1(n3850), .Y(n1642) );
  OAI22XL U2878 ( .A0(n3929), .A1(n3849), .B0(n609), .B1(n3850), .Y(n1643) );
  OAI22XL U2879 ( .A0(n3926), .A1(n3849), .B0(n610), .B1(n3850), .Y(n1644) );
  OAI22XL U2880 ( .A0(n3923), .A1(n3849), .B0(n611), .B1(n3850), .Y(n1645) );
  OAI22XL U2881 ( .A0(n3938), .A1(n3844), .B0(n639), .B1(n3845), .Y(n1673) );
  OAI22XL U2882 ( .A0(n3932), .A1(n3844), .B0(n640), .B1(n3845), .Y(n1674) );
  OAI22XL U2883 ( .A0(n3929), .A1(n175), .B0(n641), .B1(n3845), .Y(n1675) );
  OAI22XL U2884 ( .A0(n3926), .A1(n175), .B0(n642), .B1(n3845), .Y(n1676) );
  OAI22XL U2885 ( .A0(n3923), .A1(n3844), .B0(n643), .B1(n3845), .Y(n1677) );
  OAI22XL U2886 ( .A0(n3938), .A1(n3842), .B0(n671), .B1(n3843), .Y(n1705) );
  OAI22XL U2887 ( .A0(n3932), .A1(n3842), .B0(n672), .B1(n3843), .Y(n1706) );
  OAI22XL U2888 ( .A0(n3929), .A1(n3842), .B0(n673), .B1(n3843), .Y(n1707) );
  OAI22XL U2889 ( .A0(n3926), .A1(n3842), .B0(n674), .B1(n3843), .Y(n1708) );
  OAI22XL U2890 ( .A0(n3923), .A1(n3842), .B0(n675), .B1(n3843), .Y(n1709) );
  OAI22XL U2891 ( .A0(n3939), .A1(n3839), .B0(n703), .B1(n3840), .Y(n1737) );
  OAI22XL U2892 ( .A0(n3933), .A1(n3839), .B0(n704), .B1(n3840), .Y(n1738) );
  OAI22XL U2893 ( .A0(n3930), .A1(n3839), .B0(n705), .B1(n3840), .Y(n1739) );
  OAI22XL U2894 ( .A0(n3927), .A1(n3839), .B0(n706), .B1(n3840), .Y(n1740) );
  OAI22XL U2895 ( .A0(n3924), .A1(n3839), .B0(n707), .B1(n3840), .Y(n1741) );
  OAI22XL U2896 ( .A0(n3939), .A1(n3837), .B0(n735), .B1(n3838), .Y(n1769) );
  OAI22XL U2897 ( .A0(n3933), .A1(n3837), .B0(n736), .B1(n3838), .Y(n1770) );
  OAI22XL U2898 ( .A0(n3930), .A1(n3837), .B0(n737), .B1(n3838), .Y(n1771) );
  OAI22XL U2899 ( .A0(n3927), .A1(n3837), .B0(n738), .B1(n3838), .Y(n1772) );
  OAI22XL U2900 ( .A0(n3924), .A1(n3837), .B0(n739), .B1(n3838), .Y(n1773) );
  OAI22XL U2901 ( .A0(n3939), .A1(n3835), .B0(n767), .B1(n3836), .Y(n1801) );
  OAI22XL U2902 ( .A0(n3933), .A1(n3835), .B0(n768), .B1(n3836), .Y(n1802) );
  OAI22XL U2903 ( .A0(n3930), .A1(n186), .B0(n769), .B1(n3836), .Y(n1803) );
  OAI22XL U2904 ( .A0(n3927), .A1(n186), .B0(n770), .B1(n3836), .Y(n1804) );
  OAI22XL U2905 ( .A0(n3924), .A1(n3835), .B0(n771), .B1(n3836), .Y(n1805) );
  OAI22XL U2906 ( .A0(n3939), .A1(n3833), .B0(n799), .B1(n3834), .Y(n1833) );
  OAI22XL U2907 ( .A0(n3933), .A1(n3833), .B0(n800), .B1(n3834), .Y(n1834) );
  OAI22XL U2908 ( .A0(n3930), .A1(n3833), .B0(n801), .B1(n3834), .Y(n1835) );
  OAI22XL U2909 ( .A0(n3927), .A1(n3833), .B0(n802), .B1(n3834), .Y(n1836) );
  OAI22XL U2910 ( .A0(n3924), .A1(n3833), .B0(n803), .B1(n3834), .Y(n1837) );
  OAI22XL U2911 ( .A0(n3939), .A1(n3830), .B0(n831), .B1(n3831), .Y(n1865) );
  OAI22XL U2912 ( .A0(n3933), .A1(n3830), .B0(n832), .B1(n3831), .Y(n1866) );
  OAI22XL U2913 ( .A0(n3930), .A1(n191), .B0(n833), .B1(n3831), .Y(n1867) );
  OAI22XL U2914 ( .A0(n3927), .A1(n191), .B0(n834), .B1(n3831), .Y(n1868) );
  OAI22XL U2915 ( .A0(n3924), .A1(n3830), .B0(n835), .B1(n3831), .Y(n1869) );
  OAI22XL U2916 ( .A0(n3939), .A1(n3828), .B0(n863), .B1(n3829), .Y(n1897) );
  OAI22XL U2917 ( .A0(n3933), .A1(n3828), .B0(n864), .B1(n3829), .Y(n1898) );
  OAI22XL U2918 ( .A0(n3930), .A1(n3828), .B0(n865), .B1(n3829), .Y(n1899) );
  OAI22XL U2919 ( .A0(n3927), .A1(n3828), .B0(n866), .B1(n3829), .Y(n1900) );
  OAI22XL U2920 ( .A0(n3924), .A1(n3828), .B0(n867), .B1(n3829), .Y(n1901) );
  OAI22XL U2921 ( .A0(n3939), .A1(n3826), .B0(n895), .B1(n3827), .Y(n1929) );
  OAI22XL U2922 ( .A0(n3933), .A1(n3826), .B0(n896), .B1(n3827), .Y(n1930) );
  OAI22XL U2923 ( .A0(n3930), .A1(n196), .B0(n897), .B1(n3827), .Y(n1931) );
  OAI22XL U2924 ( .A0(n3927), .A1(n196), .B0(n898), .B1(n3827), .Y(n1932) );
  OAI22XL U2925 ( .A0(n3924), .A1(n3826), .B0(n899), .B1(n3827), .Y(n1933) );
  OAI22XL U2926 ( .A0(n3939), .A1(n3824), .B0(n927), .B1(n3825), .Y(n1961) );
  OAI22XL U2927 ( .A0(n3933), .A1(n3824), .B0(n928), .B1(n3825), .Y(n1962) );
  OAI22XL U2928 ( .A0(n3930), .A1(n3824), .B0(n929), .B1(n3825), .Y(n1963) );
  OAI22XL U2929 ( .A0(n3927), .A1(n3824), .B0(n930), .B1(n3825), .Y(n1964) );
  OAI22XL U2930 ( .A0(n3924), .A1(n3824), .B0(n931), .B1(n3825), .Y(n1965) );
  OAI22XL U2931 ( .A0(n3939), .A1(n3819), .B0(n959), .B1(n3820), .Y(n1993) );
  OAI22XL U2932 ( .A0(n3933), .A1(n3819), .B0(n960), .B1(n3820), .Y(n1994) );
  OAI22XL U2933 ( .A0(n3930), .A1(n204), .B0(n961), .B1(n3820), .Y(n1995) );
  OAI22XL U2934 ( .A0(n3927), .A1(n204), .B0(n962), .B1(n3820), .Y(n1996) );
  OAI22XL U2935 ( .A0(n3924), .A1(n3819), .B0(n963), .B1(n3820), .Y(n1997) );
  OAI22XL U2936 ( .A0(n3939), .A1(n3817), .B0(n991), .B1(n3818), .Y(n2025) );
  OAI22XL U2937 ( .A0(n3933), .A1(n3817), .B0(n992), .B1(n3818), .Y(n2026) );
  OAI22XL U2938 ( .A0(n3930), .A1(n3817), .B0(n993), .B1(n3818), .Y(n2027) );
  OAI22XL U2939 ( .A0(n3927), .A1(n3817), .B0(n994), .B1(n3818), .Y(n2028) );
  OAI22XL U2940 ( .A0(n3924), .A1(n3817), .B0(n995), .B1(n3818), .Y(n2029) );
  OAI22XL U2941 ( .A0(n3939), .A1(n3815), .B0(n1023), .B1(n3816), .Y(n2057) );
  OAI22XL U2942 ( .A0(n3933), .A1(n3815), .B0(n1024), .B1(n3816), .Y(n2058) );
  OAI22XL U2943 ( .A0(n3930), .A1(n209), .B0(n1025), .B1(n3816), .Y(n2059) );
  OAI22XL U2944 ( .A0(n3927), .A1(n209), .B0(n1026), .B1(n3816), .Y(n2060) );
  OAI22XL U2945 ( .A0(n3924), .A1(n3815), .B0(n1027), .B1(n3816), .Y(n2061) );
  OAI22XL U2946 ( .A0(n3940), .A1(n3813), .B0(n1055), .B1(n3814), .Y(n2089) );
  OAI22XL U2947 ( .A0(n3934), .A1(n3813), .B0(n1056), .B1(n3814), .Y(n2090) );
  OAI22XL U2948 ( .A0(n3931), .A1(n3813), .B0(n1057), .B1(n3814), .Y(n2091) );
  OAI22XL U2949 ( .A0(n3928), .A1(n3813), .B0(n1058), .B1(n3814), .Y(n2092) );
  OAI22XL U2950 ( .A0(n3925), .A1(n3813), .B0(n1059), .B1(n3814), .Y(n2093) );
  OAI22XL U2951 ( .A0(n3940), .A1(n3809), .B0(n1087), .B1(n3810), .Y(n2121) );
  OAI22XL U2952 ( .A0(n3934), .A1(n3809), .B0(n1088), .B1(n3810), .Y(n2122) );
  OAI22XL U2953 ( .A0(n3931), .A1(n214), .B0(n1089), .B1(n3810), .Y(n2123) );
  OAI22XL U2954 ( .A0(n3928), .A1(n214), .B0(n1090), .B1(n3810), .Y(n2124) );
  OAI22XL U2955 ( .A0(n3925), .A1(n3809), .B0(n1091), .B1(n3810), .Y(n2125) );
  OAI22XL U2956 ( .A0(n3940), .A1(n3806), .B0(n1119), .B1(n3807), .Y(n2153) );
  OAI22XL U2957 ( .A0(n3934), .A1(n3806), .B0(n1120), .B1(n3807), .Y(n2154) );
  OAI22XL U2958 ( .A0(n3931), .A1(n217), .B0(n1121), .B1(n3807), .Y(n2155) );
  OAI22XL U2959 ( .A0(n3928), .A1(n217), .B0(n1122), .B1(n3807), .Y(n2156) );
  OAI22XL U2960 ( .A0(n3925), .A1(n3806), .B0(n1123), .B1(n3807), .Y(n2157) );
  OAI22XL U2961 ( .A0(n3940), .A1(n3804), .B0(n1151), .B1(n3805), .Y(n2185) );
  OAI22XL U2962 ( .A0(n3934), .A1(n3804), .B0(n1152), .B1(n3805), .Y(n2186) );
  OAI22XL U2963 ( .A0(n3931), .A1(n219), .B0(n1153), .B1(n3805), .Y(n2187) );
  OAI22XL U2964 ( .A0(n3928), .A1(n219), .B0(n1154), .B1(n3805), .Y(n2188) );
  OAI22XL U2965 ( .A0(n3925), .A1(n3804), .B0(n1155), .B1(n3805), .Y(n2189) );
  OAI22XL U2966 ( .A0(n3940), .A1(n3801), .B0(n1183), .B1(n3802), .Y(n2217) );
  OAI22XL U2967 ( .A0(n3934), .A1(n3801), .B0(n1184), .B1(n3802), .Y(n2218) );
  OAI22XL U2968 ( .A0(n3931), .A1(n222), .B0(n1185), .B1(n3802), .Y(n2219) );
  OAI22XL U2969 ( .A0(n3928), .A1(n222), .B0(n1186), .B1(n3802), .Y(n2220) );
  OAI22XL U2970 ( .A0(n3925), .A1(n3801), .B0(n1187), .B1(n3802), .Y(n2221) );
  OAI22XL U2971 ( .A0(n3940), .A1(n3799), .B0(n1215), .B1(n3800), .Y(n2249) );
  OAI22XL U2972 ( .A0(n3934), .A1(n3799), .B0(n1216), .B1(n3800), .Y(n2250) );
  OAI22XL U2973 ( .A0(n3931), .A1(n225), .B0(n1217), .B1(n3800), .Y(n2251) );
  OAI22XL U2974 ( .A0(n3928), .A1(n225), .B0(n1218), .B1(n3800), .Y(n2252) );
  OAI22XL U2975 ( .A0(n3925), .A1(n3799), .B0(n1219), .B1(n3800), .Y(n2253) );
  OAI22XL U2976 ( .A0(n3938), .A1(n3962), .B0(n1279), .B1(n3963), .Y(n2313) );
  OAI22XL U2977 ( .A0(n3932), .A1(n3962), .B0(n1280), .B1(n3963), .Y(n2314) );
  OAI22XL U2978 ( .A0(n3929), .A1(n114), .B0(n1281), .B1(n3963), .Y(n2315) );
  OAI22XL U2979 ( .A0(n3926), .A1(n114), .B0(n1282), .B1(n3963), .Y(n2316) );
  OAI22XL U2980 ( .A0(n3923), .A1(n3962), .B0(n1283), .B1(n3963), .Y(n2317) );
  OAI22XL U2981 ( .A0(n3938), .A1(n3867), .B0(n1311), .B1(n3868), .Y(n2345) );
  OAI22XL U2982 ( .A0(n3932), .A1(n3867), .B0(n1312), .B1(n3868), .Y(n2346) );
  OAI22XL U2983 ( .A0(n3929), .A1(n149), .B0(n1313), .B1(n3868), .Y(n2347) );
  OAI22XL U2984 ( .A0(n3926), .A1(n149), .B0(n1314), .B1(n3868), .Y(n2348) );
  OAI22XL U2985 ( .A0(n3923), .A1(n3867), .B0(n1315), .B1(n3868), .Y(n2349) );
  OAI22XL U2986 ( .A0(n3938), .A1(n3864), .B0(n1343), .B1(n3865), .Y(n2377) );
  OAI22XL U2987 ( .A0(n3932), .A1(n3864), .B0(n1344), .B1(n3865), .Y(n2378) );
  OAI22XL U2988 ( .A0(n3929), .A1(n152), .B0(n1345), .B1(n3865), .Y(n2379) );
  OAI22XL U2989 ( .A0(n3926), .A1(n152), .B0(n1346), .B1(n3865), .Y(n2380) );
  OAI22XL U2990 ( .A0(n3923), .A1(n3864), .B0(n1347), .B1(n3865), .Y(n2381) );
  OAI22XL U2991 ( .A0(n3938), .A1(n3861), .B0(n1375), .B1(n3862), .Y(n2409) );
  OAI22XL U2992 ( .A0(n3932), .A1(n3861), .B0(n1376), .B1(n3862), .Y(n2410) );
  OAI22XL U2993 ( .A0(n3929), .A1(n156), .B0(n1377), .B1(n3862), .Y(n2411) );
  OAI22XL U2994 ( .A0(n3926), .A1(n156), .B0(n1378), .B1(n3862), .Y(n2412) );
  OAI22XL U2995 ( .A0(n3923), .A1(n3861), .B0(n1379), .B1(n3862), .Y(n2413) );
  OAI22XL U2996 ( .A0(n3938), .A1(n3858), .B0(n1407), .B1(n3859), .Y(n2441) );
  OAI22XL U2997 ( .A0(n3932), .A1(n3858), .B0(n1408), .B1(n3859), .Y(n2442) );
  OAI22XL U2998 ( .A0(n3929), .A1(n159), .B0(n1409), .B1(n3859), .Y(n2443) );
  OAI22XL U2999 ( .A0(n3926), .A1(n159), .B0(n1410), .B1(n3859), .Y(n2444) );
  OAI22XL U3000 ( .A0(n3923), .A1(n3858), .B0(n1411), .B1(n3859), .Y(n2445) );
  OAI22XL U3001 ( .A0(n3938), .A1(n3855), .B0(n1439), .B1(n3856), .Y(n2473) );
  OAI22XL U3002 ( .A0(n3932), .A1(n3855), .B0(n1440), .B1(n3856), .Y(n2474) );
  OAI22XL U3003 ( .A0(n3929), .A1(n161), .B0(n1441), .B1(n3856), .Y(n2475) );
  OAI22XL U3004 ( .A0(n3926), .A1(n161), .B0(n1442), .B1(n3856), .Y(n2476) );
  OAI22XL U3005 ( .A0(n3923), .A1(n3855), .B0(n1443), .B1(n3856), .Y(n2477) );
  OAI22XL U3006 ( .A0(n3938), .A1(n3853), .B0(n1471), .B1(n3854), .Y(n2505) );
  OAI22XL U3007 ( .A0(n3932), .A1(n3853), .B0(n1472), .B1(n3854), .Y(n2506) );
  OAI22XL U3008 ( .A0(n3929), .A1(n165), .B0(n1473), .B1(n3854), .Y(n2507) );
  OAI22XL U3009 ( .A0(n3926), .A1(n165), .B0(n1474), .B1(n3854), .Y(n2508) );
  OAI22XL U3010 ( .A0(n3923), .A1(n3853), .B0(n1475), .B1(n3854), .Y(n2509) );
  OAI22XL U3011 ( .A0(n3938), .A1(n3847), .B0(n1503), .B1(n3848), .Y(n2537) );
  OAI22XL U3012 ( .A0(n3932), .A1(n3847), .B0(n1504), .B1(n3848), .Y(n2538) );
  OAI22XL U3013 ( .A0(n3929), .A1(n3847), .B0(n1505), .B1(n3848), .Y(n2539) );
  OAI22XL U3014 ( .A0(n3926), .A1(n3847), .B0(n1506), .B1(n3848), .Y(n2540) );
  OAI22XL U3015 ( .A0(n3923), .A1(n3847), .B0(n1507), .B1(n3848), .Y(n2541) );
  OAI22XL U3016 ( .A0(n3939), .A1(n3821), .B0(n1535), .B1(n3822), .Y(n2569) );
  OAI22XL U3017 ( .A0(n3933), .A1(n3821), .B0(n1536), .B1(n3822), .Y(n2570) );
  OAI22XL U3018 ( .A0(n3930), .A1(n201), .B0(n1537), .B1(n3822), .Y(n2571) );
  OAI22XL U3019 ( .A0(n3927), .A1(n201), .B0(n1538), .B1(n3822), .Y(n2572) );
  OAI22XL U3020 ( .A0(n3924), .A1(n3821), .B0(n1539), .B1(n3822), .Y(n2573) );
  AOI222XL U3021 ( .A0(dataout[30]), .A1(n252), .B0(N958), .B1(n3776), .C0(
        n3997), .C1(n4009), .Y(n311) );
  AOI222XL U3022 ( .A0(N687), .A1(n3781), .B0(n2652), .B1(n315), .C0(N223), 
        .C1(n316), .Y(n314) );
  AOI222XL U3023 ( .A0(dataout[29]), .A1(n3772), .B0(N957), .B1(n3776), .C0(
        n3997), .C1(n2738), .Y(n325) );
  AOI222XL U3024 ( .A0(N925), .A1(n253), .B0(N893), .B1(n3778), .C0(N814), 
        .C1(n249), .Y(n326) );
  AOI222XL U3025 ( .A0(N686), .A1(n247), .B0(N192), .B1(n329), .C0(N224), .C1(
        n330), .Y(n328) );
  AOI222XL U3026 ( .A0(dataout[28]), .A1(n252), .B0(N956), .B1(n3775), .C0(
        n3997), .C1(n2696), .Y(n331) );
  AOI222XL U3027 ( .A0(N685), .A1(n3781), .B0(N193), .B1(n335), .C0(N225), 
        .C1(n336), .Y(n334) );
  AND4X1 U3028 ( .A(n337), .B(n338), .C(n339), .D(n340), .Y(n127) );
  AOI222XL U3029 ( .A0(dataout[27]), .A1(n3771), .B0(N955), .B1(n3776), .C0(
        n3997), .C1(n4010), .Y(n337) );
  AOI222XL U3030 ( .A0(N923), .A1(n253), .B0(N891), .B1(n3778), .C0(N812), 
        .C1(n249), .Y(n338) );
  AOI222XL U3031 ( .A0(N684), .A1(n247), .B0(n2651), .B1(n341), .C0(N226), 
        .C1(n342), .Y(n340) );
  AND4X1 U3032 ( .A(n343), .B(n344), .C(n345), .D(n346), .Y(n128) );
  AOI222XL U3033 ( .A0(dataout[26]), .A1(n3772), .B0(N954), .B1(n3775), .C0(
        n3997), .C1(n2704), .Y(n343) );
  AOI222XL U3034 ( .A0(N922), .A1(n3777), .B0(N890), .B1(n251), .C0(N811), 
        .C1(n3782), .Y(n344) );
  AOI222XL U3035 ( .A0(N683), .A1(n3781), .B0(N195), .B1(n347), .C0(N227), 
        .C1(n348), .Y(n346) );
  NOR2X1 U3036 ( .A(\R[3][0] ), .B(n3205), .Y(n3172) );
  NOR2X1 U3037 ( .A(\R[3][6] ), .B(n3199), .Y(n3142) );
  NOR2X1 U3038 ( .A(\R[3][5] ), .B(n3200), .Y(n3147) );
  NOR2X1 U3039 ( .A(\R[3][4] ), .B(n3201), .Y(n3152) );
  NOR2X1 U3040 ( .A(\R[3][3] ), .B(n3202), .Y(n3157) );
  NOR2X1 U3041 ( .A(\R[3][2] ), .B(n3203), .Y(n3162) );
  NOR2X1 U3042 ( .A(n3213), .B(\R[1][0] ), .Y(n3174) );
  NOR2X1 U3043 ( .A(n3213), .B(\R[1][6] ), .Y(n3144) );
  NOR2X1 U3044 ( .A(n3213), .B(\R[1][5] ), .Y(n3149) );
  NOR2X1 U3045 ( .A(n3213), .B(\R[1][4] ), .Y(n3154) );
  NOR2X1 U3046 ( .A(n3213), .B(\R[1][3] ), .Y(n3159) );
  NOR2X1 U3047 ( .A(n3213), .B(\R[1][2] ), .Y(n3164) );
  NOR2X1 U3048 ( .A(n3213), .B(\R[1][1] ), .Y(n3169) );
  MXI4X1 U3049 ( .A(n3271), .B(n3272), .C(n3273), .D(n3274), .S0(n3760), .S1(
        n3752), .Y(n3270) );
  MXI4X1 U3050 ( .A(n3266), .B(n3267), .C(n3268), .D(n3269), .S0(n3760), .S1(
        n3752), .Y(n3265) );
  CLKMX2X2 U3051 ( .A(n3260), .B(n3255), .S0(n3767), .Y(N251) );
  MXI4X1 U3052 ( .A(n3261), .B(n3262), .C(n3263), .D(n3264), .S0(n3760), .S1(
        n3752), .Y(n3260) );
  MXI4X1 U3053 ( .A(n3256), .B(n3257), .C(n3258), .D(n3259), .S0(n3760), .S1(
        n3752), .Y(n3255) );
  MXI4X1 U3054 ( .A(\R[12][2] ), .B(\R[13][2] ), .C(\R[14][2] ), .D(\R[15][2] ), .S0(n3717), .S1(n3742), .Y(n3264) );
  CLKMX2X2 U3055 ( .A(n3250), .B(n3245), .S0(n3767), .Y(N252) );
  MXI4X1 U3056 ( .A(n3251), .B(n3252), .C(n3253), .D(n3254), .S0(n3759), .S1(
        n3751), .Y(n3250) );
  MXI4X1 U3057 ( .A(n3246), .B(n3247), .C(n3248), .D(n3249), .S0(n3759), .S1(
        n3751), .Y(n3245) );
  MXI4X1 U3058 ( .A(\R[12][1] ), .B(\R[13][1] ), .C(\R[14][1] ), .D(\R[15][1] ), .S0(n3717), .S1(n3742), .Y(n3254) );
  CLKMX2X2 U3059 ( .A(n3240), .B(n3235), .S0(n3767), .Y(N253) );
  MXI4X1 U3060 ( .A(n3236), .B(n3237), .C(n3238), .D(n3239), .S0(n3759), .S1(
        n3751), .Y(n3235) );
  MXI4X1 U3061 ( .A(n3241), .B(n3242), .C(n3243), .D(n3244), .S0(n3759), .S1(
        n3751), .Y(n3240) );
  MXI4X1 U3062 ( .A(\R[28][0] ), .B(\R[29][0] ), .C(\R[30][0] ), .D(\R[31][0] ), .S0(n3717), .S1(n3742), .Y(n3239) );
  MXI4X1 U3063 ( .A(\R[20][0] ), .B(\R[21][0] ), .C(\R[22][0] ), .D(\R[23][0] ), .S0(n3179), .S1(n3206), .Y(n2763) );
  MXI4X1 U3064 ( .A(\R[4][0] ), .B(\R[5][0] ), .C(\R[6][0] ), .D(\R[7][0] ), 
        .S0(n3179), .S1(n3206), .Y(n2767) );
  MXI4X1 U3065 ( .A(\R[20][6] ), .B(\R[21][6] ), .C(\R[22][6] ), .D(\R[23][6] ), .S0(n3180), .S1(n3207), .Y(n2811) );
  MXI4X1 U3066 ( .A(\R[4][6] ), .B(\R[5][6] ), .C(\R[6][6] ), .D(\R[7][6] ), 
        .S0(n3180), .S1(n3207), .Y(n2815) );
  MXI4X1 U3067 ( .A(\R[4][5] ), .B(\R[5][5] ), .C(\R[6][5] ), .D(\R[7][5] ), 
        .S0(n3180), .S1(n3207), .Y(n2807) );
  MXI4X1 U3068 ( .A(\R[20][4] ), .B(\R[21][4] ), .C(\R[22][4] ), .D(\R[23][4] ), .S0(n3179), .S1(n3207), .Y(n2795) );
  MXI4X1 U3069 ( .A(\R[4][4] ), .B(\R[5][4] ), .C(\R[6][4] ), .D(\R[7][4] ), 
        .S0(n3179), .S1(n3207), .Y(n2799) );
  MXI4X1 U3070 ( .A(\R[20][3] ), .B(\R[21][3] ), .C(\R[22][3] ), .D(\R[23][3] ), .S0(n3179), .S1(n3206), .Y(n2787) );
  MXI4X1 U3071 ( .A(\R[4][3] ), .B(\R[5][3] ), .C(\R[6][3] ), .D(\R[7][3] ), 
        .S0(n3179), .S1(n3206), .Y(n2791) );
  MXI4X1 U3072 ( .A(\R[20][2] ), .B(\R[21][2] ), .C(\R[22][2] ), .D(\R[23][2] ), .S0(n3179), .S1(n3206), .Y(n2779) );
  MXI4X1 U3073 ( .A(\R[4][2] ), .B(\R[5][2] ), .C(\R[6][2] ), .D(\R[7][2] ), 
        .S0(n3179), .S1(n3206), .Y(n2783) );
  MXI4X1 U3074 ( .A(\R[16][0] ), .B(\R[17][0] ), .C(\R[18][0] ), .D(\R[19][0] ), .S0(n3179), .S1(n3206), .Y(n2761) );
  MXI4X1 U3075 ( .A(\R[16][6] ), .B(\R[17][6] ), .C(\R[18][6] ), .D(\R[19][6] ), .S0(n3180), .S1(n3207), .Y(n2809) );
  MXI4X1 U3076 ( .A(\R[16][4] ), .B(\R[17][4] ), .C(\R[18][4] ), .D(\R[19][4] ), .S0(n3179), .S1(n3207), .Y(n2793) );
  MXI4X1 U3077 ( .A(\R[16][3] ), .B(\R[17][3] ), .C(\R[18][3] ), .D(\R[19][3] ), .S0(n3179), .S1(n3206), .Y(n2785) );
  MXI4X1 U3078 ( .A(\R[16][2] ), .B(\R[17][2] ), .C(\R[18][2] ), .D(\R[19][2] ), .S0(n3179), .S1(n3206), .Y(n2777) );
  MXI4X1 U3079 ( .A(\R[24][0] ), .B(\R[25][0] ), .C(\R[26][0] ), .D(\R[27][0] ), .S0(n3179), .S1(n3206), .Y(n2762) );
  MXI4X1 U3080 ( .A(\R[8][0] ), .B(\R[9][0] ), .C(\R[10][0] ), .D(\R[11][0] ), 
        .S0(n3179), .S1(n3206), .Y(n2766) );
  MXI4X1 U3081 ( .A(\R[24][6] ), .B(\R[25][6] ), .C(\R[26][6] ), .D(\R[27][6] ), .S0(n3180), .S1(n3207), .Y(n2810) );
  MXI4X1 U3082 ( .A(\R[8][6] ), .B(\R[9][6] ), .C(\R[10][6] ), .D(\R[11][6] ), 
        .S0(n3180), .S1(n3207), .Y(n2814) );
  MXI4X1 U3083 ( .A(\R[8][5] ), .B(\R[9][5] ), .C(\R[10][5] ), .D(\R[11][5] ), 
        .S0(n3180), .S1(n3207), .Y(n2806) );
  MXI4X1 U3084 ( .A(\R[24][3] ), .B(\R[25][3] ), .C(\R[26][3] ), .D(\R[27][3] ), .S0(n3179), .S1(n3206), .Y(n2786) );
  MXI4X1 U3085 ( .A(\R[8][3] ), .B(\R[9][3] ), .C(\R[10][3] ), .D(\R[11][3] ), 
        .S0(n3179), .S1(n3206), .Y(n2790) );
  MXI4X1 U3086 ( .A(\R[24][2] ), .B(\R[25][2] ), .C(\R[26][2] ), .D(\R[27][2] ), .S0(n3179), .S1(n3206), .Y(n2778) );
  MXI4X1 U3087 ( .A(\R[8][2] ), .B(\R[9][2] ), .C(\R[10][2] ), .D(\R[11][2] ), 
        .S0(n3179), .S1(n3206), .Y(n2782) );
  MXI4X1 U3088 ( .A(\R[28][0] ), .B(\R[29][0] ), .C(\R[30][0] ), .D(\R[31][0] ), .S0(n3179), .S1(n3206), .Y(n2764) );
  MXI4X1 U3089 ( .A(\R[12][0] ), .B(\R[13][0] ), .C(\R[14][0] ), .D(\R[15][0] ), .S0(n3179), .S1(n3206), .Y(n2768) );
  MXI4X1 U3090 ( .A(\R[28][6] ), .B(\R[29][6] ), .C(\R[30][6] ), .D(\R[31][6] ), .S0(n3180), .S1(n3207), .Y(n2812) );
  MXI4X1 U3091 ( .A(\R[12][6] ), .B(\R[13][6] ), .C(\R[14][6] ), .D(\R[15][6] ), .S0(n3180), .S1(n3207), .Y(n2816) );
  MXI4X1 U3092 ( .A(\R[28][4] ), .B(\R[29][4] ), .C(\R[30][4] ), .D(\R[31][4] ), .S0(n3179), .S1(n3207), .Y(n2796) );
  MXI4X1 U3093 ( .A(\R[12][4] ), .B(\R[13][4] ), .C(\R[14][4] ), .D(\R[15][4] ), .S0(n3179), .S1(n3207), .Y(n2800) );
  MXI4X1 U3094 ( .A(\R[28][3] ), .B(\R[29][3] ), .C(\R[30][3] ), .D(\R[31][3] ), .S0(n3179), .S1(n3206), .Y(n2788) );
  MXI4X1 U3095 ( .A(\R[12][3] ), .B(\R[13][3] ), .C(\R[14][3] ), .D(\R[15][3] ), .S0(n3179), .S1(n3206), .Y(n2792) );
  MXI4X1 U3096 ( .A(\R[28][2] ), .B(\R[29][2] ), .C(\R[30][2] ), .D(\R[31][2] ), .S0(n3179), .S1(n3206), .Y(n2780) );
  MXI4X1 U3097 ( .A(\R[12][2] ), .B(\R[13][2] ), .C(\R[14][2] ), .D(\R[15][2] ), .S0(n3179), .S1(n3206), .Y(n2784) );
  MXI4X1 U3098 ( .A(\R[12][1] ), .B(\R[13][1] ), .C(\R[14][1] ), .D(\R[15][1] ), .S0(n3179), .S1(n3206), .Y(n2776) );
  CLKMX2X2 U3099 ( .A(n3310), .B(n3305), .S0(n3767), .Y(N246) );
  MXI4X1 U3100 ( .A(n3311), .B(n3312), .C(n3313), .D(n3314), .S0(n3760), .S1(
        n3752), .Y(n3310) );
  MXI4X1 U3101 ( .A(n3306), .B(n3307), .C(n3308), .D(n3309), .S0(n3760), .S1(
        n3752), .Y(n3305) );
  MXI4X1 U3102 ( .A(\R[12][7] ), .B(\R[13][7] ), .C(\R[14][7] ), .D(\R[15][7] ), .S0(n3718), .S1(n3743), .Y(n3314) );
  CLKMX2X2 U3103 ( .A(n3300), .B(n3295), .S0(n3767), .Y(N247) );
  MXI4X1 U3104 ( .A(n3301), .B(n3302), .C(n3303), .D(n3304), .S0(n3760), .S1(
        n3752), .Y(n3300) );
  MXI4X1 U3105 ( .A(n3296), .B(n3297), .C(n3298), .D(n3299), .S0(n3760), .S1(
        n3752), .Y(n3295) );
  MXI4X1 U3106 ( .A(\R[12][6] ), .B(\R[13][6] ), .C(\R[14][6] ), .D(\R[15][6] ), .S0(n3718), .S1(n3743), .Y(n3304) );
  CLKMX2X2 U3107 ( .A(n3340), .B(n3335), .S0(n3768), .Y(N243) );
  MXI4X1 U3108 ( .A(n3341), .B(n3342), .C(n3343), .D(n3344), .S0(n3761), .S1(
        n3753), .Y(n3340) );
  MXI4X1 U3109 ( .A(n3336), .B(n3337), .C(n3338), .D(n3339), .S0(n3761), .S1(
        n3753), .Y(n3335) );
  MXI4X1 U3110 ( .A(\R[12][10] ), .B(\R[13][10] ), .C(\R[14][10] ), .D(
        \R[15][10] ), .S0(n3718), .S1(n3743), .Y(n3344) );
  CLKMX2X2 U3111 ( .A(n3320), .B(n3315), .S0(n3768), .Y(N245) );
  MXI4X1 U3112 ( .A(n3321), .B(n3322), .C(n3323), .D(n3324), .S0(n3761), .S1(
        n3753), .Y(n3320) );
  MXI4X1 U3113 ( .A(n3316), .B(n3317), .C(n3318), .D(n3319), .S0(n3761), .S1(
        n3753), .Y(n3315) );
  MXI4X1 U3114 ( .A(\R[12][8] ), .B(\R[13][8] ), .C(\R[14][8] ), .D(\R[15][8] ), .S0(n3718), .S1(n3743), .Y(n3324) );
  CLKMX2X2 U3115 ( .A(n3350), .B(n3345), .S0(n3768), .Y(N242) );
  MXI4X1 U3116 ( .A(n3351), .B(n3352), .C(n3353), .D(n3354), .S0(n3761), .S1(
        n3753), .Y(n3350) );
  MXI4X1 U3117 ( .A(n3346), .B(n3347), .C(n3348), .D(n3349), .S0(n3761), .S1(
        n3753), .Y(n3345) );
  MXI4X1 U3118 ( .A(\R[12][11] ), .B(\R[13][11] ), .C(\R[14][11] ), .D(
        \R[15][11] ), .S0(n3718), .S1(n3743), .Y(n3354) );
  CLKMX2X2 U3119 ( .A(n3330), .B(n3325), .S0(n3768), .Y(N244) );
  MXI4X1 U3120 ( .A(n3331), .B(n3332), .C(n3333), .D(n3334), .S0(n3761), .S1(
        n3753), .Y(n3330) );
  MXI4X1 U3121 ( .A(n3326), .B(n3327), .C(n3328), .D(n3329), .S0(n3761), .S1(
        n3753), .Y(n3325) );
  MXI4X1 U3122 ( .A(\R[12][9] ), .B(\R[13][9] ), .C(\R[14][9] ), .D(\R[15][9] ), .S0(n3718), .S1(n3743), .Y(n3334) );
  NOR2X1 U3123 ( .A(instruction[28]), .B(instruction[29]), .Y(n552) );
  OAI22XL U3124 ( .A0(n3920), .A1(n3851), .B0(n580), .B1(n3852), .Y(n1614) );
  OAI22XL U3125 ( .A0(n3917), .A1(n3851), .B0(n581), .B1(n3852), .Y(n1615) );
  OAI22XL U3126 ( .A0(n3914), .A1(n3851), .B0(n582), .B1(n3852), .Y(n1616) );
  OAI22XL U3127 ( .A0(n3911), .A1(n3851), .B0(n583), .B1(n3852), .Y(n1617) );
  OAI22XL U3128 ( .A0(n3908), .A1(n3851), .B0(n584), .B1(n3852), .Y(n1618) );
  OAI22XL U3129 ( .A0(n3905), .A1(n3851), .B0(n585), .B1(n3852), .Y(n1619) );
  OAI22XL U3130 ( .A0(n3920), .A1(n3849), .B0(n612), .B1(n3850), .Y(n1646) );
  OAI22XL U3131 ( .A0(n3917), .A1(n3849), .B0(n613), .B1(n3850), .Y(n1647) );
  OAI22XL U3132 ( .A0(n3914), .A1(n3849), .B0(n614), .B1(n3850), .Y(n1648) );
  OAI22XL U3133 ( .A0(n3911), .A1(n3849), .B0(n615), .B1(n3850), .Y(n1649) );
  OAI22XL U3134 ( .A0(n3908), .A1(n3849), .B0(n616), .B1(n3850), .Y(n1650) );
  OAI22XL U3135 ( .A0(n3905), .A1(n3849), .B0(n617), .B1(n3850), .Y(n1651) );
  OAI22XL U3136 ( .A0(n3920), .A1(n3844), .B0(n644), .B1(n3845), .Y(n1678) );
  OAI22XL U3137 ( .A0(n3917), .A1(n3844), .B0(n645), .B1(n3845), .Y(n1679) );
  OAI22XL U3138 ( .A0(n3914), .A1(n3844), .B0(n646), .B1(n3845), .Y(n1680) );
  OAI22XL U3139 ( .A0(n3911), .A1(n3844), .B0(n647), .B1(n3845), .Y(n1681) );
  OAI22XL U3140 ( .A0(n3908), .A1(n3844), .B0(n648), .B1(n3845), .Y(n1682) );
  OAI22XL U3141 ( .A0(n3905), .A1(n3844), .B0(n649), .B1(n3845), .Y(n1683) );
  OAI22XL U3142 ( .A0(n3920), .A1(n3842), .B0(n676), .B1(n3843), .Y(n1710) );
  OAI22XL U3143 ( .A0(n3917), .A1(n3842), .B0(n677), .B1(n3843), .Y(n1711) );
  OAI22XL U3144 ( .A0(n3914), .A1(n3842), .B0(n678), .B1(n3843), .Y(n1712) );
  OAI22XL U3145 ( .A0(n3911), .A1(n3842), .B0(n679), .B1(n3843), .Y(n1713) );
  OAI22XL U3146 ( .A0(n3908), .A1(n3842), .B0(n680), .B1(n3843), .Y(n1714) );
  OAI22XL U3147 ( .A0(n3905), .A1(n3841), .B0(n681), .B1(n3843), .Y(n1715) );
  OAI22XL U3148 ( .A0(n3921), .A1(n3839), .B0(n708), .B1(n3840), .Y(n1742) );
  OAI22XL U3149 ( .A0(n3918), .A1(n3839), .B0(n709), .B1(n3840), .Y(n1743) );
  OAI22XL U3150 ( .A0(n3915), .A1(n3839), .B0(n710), .B1(n3840), .Y(n1744) );
  OAI22XL U3151 ( .A0(n3912), .A1(n3839), .B0(n711), .B1(n3840), .Y(n1745) );
  OAI22XL U3152 ( .A0(n3909), .A1(n3839), .B0(n712), .B1(n3840), .Y(n1746) );
  OAI22XL U3153 ( .A0(n3906), .A1(n3839), .B0(n713), .B1(n3840), .Y(n1747) );
  OAI22XL U3154 ( .A0(n3921), .A1(n3837), .B0(n740), .B1(n3838), .Y(n1774) );
  OAI22XL U3155 ( .A0(n3918), .A1(n3837), .B0(n741), .B1(n3838), .Y(n1775) );
  OAI22XL U3156 ( .A0(n3915), .A1(n3837), .B0(n742), .B1(n3838), .Y(n1776) );
  OAI22XL U3157 ( .A0(n3912), .A1(n3837), .B0(n743), .B1(n3838), .Y(n1777) );
  OAI22XL U3158 ( .A0(n3909), .A1(n3837), .B0(n744), .B1(n3838), .Y(n1778) );
  OAI22XL U3159 ( .A0(n3906), .A1(n3837), .B0(n745), .B1(n3838), .Y(n1779) );
  OAI22XL U3160 ( .A0(n3921), .A1(n3835), .B0(n772), .B1(n3836), .Y(n1806) );
  OAI22XL U3161 ( .A0(n3918), .A1(n3835), .B0(n773), .B1(n3836), .Y(n1807) );
  OAI22XL U3162 ( .A0(n3915), .A1(n3835), .B0(n774), .B1(n3836), .Y(n1808) );
  OAI22XL U3163 ( .A0(n3912), .A1(n3835), .B0(n775), .B1(n3836), .Y(n1809) );
  OAI22XL U3164 ( .A0(n3909), .A1(n3835), .B0(n776), .B1(n3836), .Y(n1810) );
  OAI22XL U3165 ( .A0(n3906), .A1(n3835), .B0(n777), .B1(n3836), .Y(n1811) );
  OAI22XL U3166 ( .A0(n3921), .A1(n3833), .B0(n804), .B1(n3834), .Y(n1838) );
  OAI22XL U3167 ( .A0(n3918), .A1(n3833), .B0(n805), .B1(n3834), .Y(n1839) );
  OAI22XL U3168 ( .A0(n3915), .A1(n3833), .B0(n806), .B1(n3834), .Y(n1840) );
  OAI22XL U3169 ( .A0(n3912), .A1(n3833), .B0(n807), .B1(n3834), .Y(n1841) );
  OAI22XL U3170 ( .A0(n3909), .A1(n3833), .B0(n808), .B1(n3834), .Y(n1842) );
  OAI22XL U3171 ( .A0(n3906), .A1(n3832), .B0(n809), .B1(n3834), .Y(n1843) );
  OAI22XL U3172 ( .A0(n3921), .A1(n3830), .B0(n836), .B1(n3831), .Y(n1870) );
  OAI22XL U3173 ( .A0(n3918), .A1(n3830), .B0(n837), .B1(n3831), .Y(n1871) );
  OAI22XL U3174 ( .A0(n3915), .A1(n3830), .B0(n838), .B1(n3831), .Y(n1872) );
  OAI22XL U3175 ( .A0(n3912), .A1(n3830), .B0(n839), .B1(n3831), .Y(n1873) );
  OAI22XL U3176 ( .A0(n3909), .A1(n3830), .B0(n840), .B1(n3831), .Y(n1874) );
  OAI22XL U3177 ( .A0(n3906), .A1(n3830), .B0(n841), .B1(n3831), .Y(n1875) );
  OAI22XL U3178 ( .A0(n3921), .A1(n3828), .B0(n868), .B1(n3829), .Y(n1902) );
  OAI22XL U3179 ( .A0(n3918), .A1(n3828), .B0(n869), .B1(n3829), .Y(n1903) );
  OAI22XL U3180 ( .A0(n3915), .A1(n3828), .B0(n870), .B1(n3829), .Y(n1904) );
  OAI22XL U3181 ( .A0(n3912), .A1(n3828), .B0(n871), .B1(n3829), .Y(n1905) );
  OAI22XL U3182 ( .A0(n3909), .A1(n3828), .B0(n872), .B1(n3829), .Y(n1906) );
  OAI22XL U3183 ( .A0(n3906), .A1(n3828), .B0(n873), .B1(n3829), .Y(n1907) );
  OAI22XL U3184 ( .A0(n3921), .A1(n3826), .B0(n900), .B1(n3827), .Y(n1934) );
  OAI22XL U3185 ( .A0(n3918), .A1(n3826), .B0(n901), .B1(n3827), .Y(n1935) );
  OAI22XL U3186 ( .A0(n3915), .A1(n3826), .B0(n902), .B1(n3827), .Y(n1936) );
  OAI22XL U3187 ( .A0(n3912), .A1(n3826), .B0(n903), .B1(n3827), .Y(n1937) );
  OAI22XL U3188 ( .A0(n3909), .A1(n3826), .B0(n904), .B1(n3827), .Y(n1938) );
  OAI22XL U3189 ( .A0(n3906), .A1(n3826), .B0(n905), .B1(n3827), .Y(n1939) );
  OAI22XL U3190 ( .A0(n3921), .A1(n3824), .B0(n932), .B1(n3825), .Y(n1966) );
  OAI22XL U3191 ( .A0(n3918), .A1(n3824), .B0(n933), .B1(n3825), .Y(n1967) );
  OAI22XL U3192 ( .A0(n3915), .A1(n3824), .B0(n934), .B1(n3825), .Y(n1968) );
  OAI22XL U3193 ( .A0(n3912), .A1(n3824), .B0(n935), .B1(n3825), .Y(n1969) );
  OAI22XL U3194 ( .A0(n3909), .A1(n3824), .B0(n936), .B1(n3825), .Y(n1970) );
  OAI22XL U3195 ( .A0(n3906), .A1(n3823), .B0(n937), .B1(n3825), .Y(n1971) );
  OAI22XL U3196 ( .A0(n3921), .A1(n3819), .B0(n964), .B1(n3820), .Y(n1998) );
  OAI22XL U3197 ( .A0(n3918), .A1(n3819), .B0(n965), .B1(n3820), .Y(n1999) );
  OAI22XL U3198 ( .A0(n3915), .A1(n3819), .B0(n966), .B1(n3820), .Y(n2000) );
  OAI22XL U3199 ( .A0(n3912), .A1(n3819), .B0(n967), .B1(n3820), .Y(n2001) );
  OAI22XL U3200 ( .A0(n3909), .A1(n3819), .B0(n968), .B1(n3820), .Y(n2002) );
  OAI22XL U3201 ( .A0(n3906), .A1(n3819), .B0(n969), .B1(n3820), .Y(n2003) );
  OAI22XL U3202 ( .A0(n3921), .A1(n3817), .B0(n996), .B1(n3818), .Y(n2030) );
  OAI22XL U3203 ( .A0(n3918), .A1(n3817), .B0(n997), .B1(n3818), .Y(n2031) );
  OAI22XL U3204 ( .A0(n3915), .A1(n3817), .B0(n998), .B1(n3818), .Y(n2032) );
  OAI22XL U3205 ( .A0(n3912), .A1(n3817), .B0(n999), .B1(n3818), .Y(n2033) );
  OAI22XL U3206 ( .A0(n3909), .A1(n3817), .B0(n1000), .B1(n3818), .Y(n2034) );
  OAI22XL U3207 ( .A0(n3906), .A1(n3817), .B0(n1001), .B1(n3818), .Y(n2035) );
  OAI22XL U3208 ( .A0(n3921), .A1(n3815), .B0(n1028), .B1(n3816), .Y(n2062) );
  OAI22XL U3209 ( .A0(n3918), .A1(n3815), .B0(n1029), .B1(n3816), .Y(n2063) );
  OAI22XL U3210 ( .A0(n3915), .A1(n3815), .B0(n1030), .B1(n3816), .Y(n2064) );
  OAI22XL U3211 ( .A0(n3912), .A1(n3815), .B0(n1031), .B1(n3816), .Y(n2065) );
  OAI22XL U3212 ( .A0(n3909), .A1(n3815), .B0(n1032), .B1(n3816), .Y(n2066) );
  OAI22XL U3213 ( .A0(n3906), .A1(n3815), .B0(n1033), .B1(n3816), .Y(n2067) );
  OAI22XL U3214 ( .A0(n3922), .A1(n3813), .B0(n1060), .B1(n3814), .Y(n2094) );
  OAI22XL U3215 ( .A0(n3919), .A1(n3813), .B0(n1061), .B1(n3814), .Y(n2095) );
  OAI22XL U3216 ( .A0(n3916), .A1(n3813), .B0(n1062), .B1(n3814), .Y(n2096) );
  OAI22XL U3217 ( .A0(n3913), .A1(n3813), .B0(n1063), .B1(n3814), .Y(n2097) );
  OAI22XL U3218 ( .A0(n3910), .A1(n3813), .B0(n1064), .B1(n3814), .Y(n2098) );
  OAI22XL U3219 ( .A0(n3907), .A1(n3812), .B0(n1065), .B1(n3814), .Y(n2099) );
  OAI22XL U3220 ( .A0(n3922), .A1(n3809), .B0(n1092), .B1(n3810), .Y(n2126) );
  OAI22XL U3221 ( .A0(n3919), .A1(n3809), .B0(n1093), .B1(n3810), .Y(n2127) );
  OAI22XL U3222 ( .A0(n3916), .A1(n3809), .B0(n1094), .B1(n3810), .Y(n2128) );
  OAI22XL U3223 ( .A0(n3913), .A1(n3809), .B0(n1095), .B1(n3810), .Y(n2129) );
  OAI22XL U3224 ( .A0(n3910), .A1(n214), .B0(n1096), .B1(n3810), .Y(n2130) );
  OAI22XL U3225 ( .A0(n3907), .A1(n214), .B0(n1097), .B1(n3811), .Y(n2131) );
  OAI22XL U3226 ( .A0(n3922), .A1(n3806), .B0(n1124), .B1(n3807), .Y(n2158) );
  OAI22XL U3227 ( .A0(n3919), .A1(n3806), .B0(n1125), .B1(n3807), .Y(n2159) );
  OAI22XL U3228 ( .A0(n3916), .A1(n3806), .B0(n1126), .B1(n3807), .Y(n2160) );
  OAI22XL U3229 ( .A0(n3913), .A1(n3806), .B0(n1127), .B1(n3807), .Y(n2161) );
  OAI22XL U3230 ( .A0(n3910), .A1(n217), .B0(n1128), .B1(n3807), .Y(n2162) );
  OAI22XL U3231 ( .A0(n3907), .A1(n217), .B0(n1129), .B1(n3808), .Y(n2163) );
  OAI22XL U3232 ( .A0(n3922), .A1(n3804), .B0(n1156), .B1(n3805), .Y(n2190) );
  OAI22XL U3233 ( .A0(n3919), .A1(n3804), .B0(n1157), .B1(n3805), .Y(n2191) );
  OAI22XL U3234 ( .A0(n3916), .A1(n3804), .B0(n1158), .B1(n3805), .Y(n2192) );
  OAI22XL U3235 ( .A0(n3913), .A1(n3804), .B0(n1159), .B1(n3805), .Y(n2193) );
  OAI22XL U3236 ( .A0(n3910), .A1(n219), .B0(n1160), .B1(n3805), .Y(n2194) );
  OAI22XL U3237 ( .A0(n3907), .A1(n219), .B0(n1161), .B1(n3805), .Y(n2195) );
  OAI22XL U3238 ( .A0(n3922), .A1(n3801), .B0(n1188), .B1(n3802), .Y(n2222) );
  OAI22XL U3239 ( .A0(n3919), .A1(n3801), .B0(n1189), .B1(n3802), .Y(n2223) );
  OAI22XL U3240 ( .A0(n3916), .A1(n3801), .B0(n1190), .B1(n3802), .Y(n2224) );
  OAI22XL U3241 ( .A0(n3913), .A1(n3801), .B0(n1191), .B1(n3802), .Y(n2225) );
  OAI22XL U3242 ( .A0(n3910), .A1(n222), .B0(n1192), .B1(n3802), .Y(n2226) );
  OAI22XL U3243 ( .A0(n3907), .A1(n222), .B0(n1193), .B1(n3803), .Y(n2227) );
  OAI22XL U3244 ( .A0(n3922), .A1(n3799), .B0(n1220), .B1(n3800), .Y(n2254) );
  OAI22XL U3245 ( .A0(n3919), .A1(n3799), .B0(n1221), .B1(n3800), .Y(n2255) );
  OAI22XL U3246 ( .A0(n3916), .A1(n3799), .B0(n1222), .B1(n3800), .Y(n2256) );
  OAI22XL U3247 ( .A0(n3913), .A1(n3799), .B0(n1223), .B1(n3800), .Y(n2257) );
  OAI22XL U3248 ( .A0(n3910), .A1(n225), .B0(n1224), .B1(n3800), .Y(n2258) );
  OAI22XL U3249 ( .A0(n3907), .A1(n225), .B0(n1225), .B1(n3800), .Y(n2259) );
  OAI22XL U3250 ( .A0(n1253), .A1(n3798), .B0(n3919), .B1(n3796), .Y(n2287) );
  OAI22XL U3251 ( .A0(n1254), .A1(n3798), .B0(n3916), .B1(n3796), .Y(n2288) );
  OAI22XL U3252 ( .A0(n1255), .A1(n3798), .B0(n3913), .B1(n3796), .Y(n2289) );
  OAI22XL U3253 ( .A0(n1256), .A1(n3798), .B0(n3910), .B1(n3796), .Y(n2290) );
  OAI22XL U3254 ( .A0(n1257), .A1(n3798), .B0(n3907), .B1(n3797), .Y(n2291) );
  OAI22XL U3255 ( .A0(n3920), .A1(n3962), .B0(n1284), .B1(n3963), .Y(n2318) );
  OAI22XL U3256 ( .A0(n3917), .A1(n3962), .B0(n1285), .B1(n3963), .Y(n2319) );
  OAI22XL U3257 ( .A0(n3914), .A1(n3962), .B0(n1286), .B1(n3963), .Y(n2320) );
  OAI22XL U3258 ( .A0(n3911), .A1(n3962), .B0(n1287), .B1(n3963), .Y(n2321) );
  OAI22XL U3259 ( .A0(n3908), .A1(n114), .B0(n1288), .B1(n3963), .Y(n2322) );
  OAI22XL U3260 ( .A0(n3905), .A1(n114), .B0(n1289), .B1(n3963), .Y(n2323) );
  OAI22XL U3261 ( .A0(n3920), .A1(n3867), .B0(n1316), .B1(n3868), .Y(n2350) );
  OAI22XL U3262 ( .A0(n3917), .A1(n3867), .B0(n1317), .B1(n3868), .Y(n2351) );
  OAI22XL U3263 ( .A0(n3914), .A1(n3867), .B0(n1318), .B1(n3868), .Y(n2352) );
  OAI22XL U3264 ( .A0(n3911), .A1(n3867), .B0(n1319), .B1(n3868), .Y(n2353) );
  OAI22XL U3265 ( .A0(n3908), .A1(n149), .B0(n1320), .B1(n3868), .Y(n2354) );
  OAI22XL U3266 ( .A0(n3905), .A1(n149), .B0(n1321), .B1(n3868), .Y(n2355) );
  OAI22XL U3267 ( .A0(n3920), .A1(n3864), .B0(n1348), .B1(n3865), .Y(n2382) );
  OAI22XL U3268 ( .A0(n3917), .A1(n3864), .B0(n1349), .B1(n3865), .Y(n2383) );
  OAI22XL U3269 ( .A0(n3914), .A1(n3864), .B0(n1350), .B1(n3865), .Y(n2384) );
  OAI22XL U3270 ( .A0(n3911), .A1(n3864), .B0(n1351), .B1(n3865), .Y(n2385) );
  OAI22XL U3271 ( .A0(n3908), .A1(n152), .B0(n1352), .B1(n3865), .Y(n2386) );
  OAI22XL U3272 ( .A0(n3905), .A1(n152), .B0(n1353), .B1(n3866), .Y(n2387) );
  OAI22XL U3273 ( .A0(n3920), .A1(n3861), .B0(n1380), .B1(n3862), .Y(n2414) );
  OAI22XL U3274 ( .A0(n3917), .A1(n3861), .B0(n1381), .B1(n3862), .Y(n2415) );
  OAI22XL U3275 ( .A0(n3914), .A1(n3861), .B0(n1382), .B1(n3862), .Y(n2416) );
  OAI22XL U3276 ( .A0(n3911), .A1(n3861), .B0(n1383), .B1(n3862), .Y(n2417) );
  OAI22XL U3277 ( .A0(n3908), .A1(n156), .B0(n1384), .B1(n3862), .Y(n2418) );
  OAI22XL U3278 ( .A0(n3905), .A1(n156), .B0(n1385), .B1(n3863), .Y(n2419) );
  OAI22XL U3279 ( .A0(n3920), .A1(n3858), .B0(n1412), .B1(n3859), .Y(n2446) );
  OAI22XL U3280 ( .A0(n3917), .A1(n3858), .B0(n1413), .B1(n3859), .Y(n2447) );
  OAI22XL U3281 ( .A0(n3914), .A1(n3858), .B0(n1414), .B1(n3859), .Y(n2448) );
  OAI22XL U3282 ( .A0(n3911), .A1(n3858), .B0(n1415), .B1(n3859), .Y(n2449) );
  OAI22XL U3283 ( .A0(n3908), .A1(n159), .B0(n1416), .B1(n3859), .Y(n2450) );
  OAI22XL U3284 ( .A0(n3905), .A1(n159), .B0(n1417), .B1(n3860), .Y(n2451) );
  OAI22XL U3285 ( .A0(n3920), .A1(n3855), .B0(n1444), .B1(n3856), .Y(n2478) );
  OAI22XL U3286 ( .A0(n3917), .A1(n3855), .B0(n1445), .B1(n3856), .Y(n2479) );
  OAI22XL U3287 ( .A0(n3914), .A1(n3855), .B0(n1446), .B1(n3856), .Y(n2480) );
  OAI22XL U3288 ( .A0(n3911), .A1(n3855), .B0(n1447), .B1(n3856), .Y(n2481) );
  OAI22XL U3289 ( .A0(n3908), .A1(n161), .B0(n1448), .B1(n3856), .Y(n2482) );
  OAI22XL U3290 ( .A0(n3905), .A1(n161), .B0(n1449), .B1(n3857), .Y(n2483) );
  OAI22XL U3291 ( .A0(n3920), .A1(n3853), .B0(n1476), .B1(n3854), .Y(n2510) );
  OAI22XL U3292 ( .A0(n3917), .A1(n3853), .B0(n1477), .B1(n3854), .Y(n2511) );
  OAI22XL U3293 ( .A0(n3914), .A1(n3853), .B0(n1478), .B1(n3854), .Y(n2512) );
  OAI22XL U3294 ( .A0(n3911), .A1(n3853), .B0(n1479), .B1(n3854), .Y(n2513) );
  OAI22XL U3295 ( .A0(n3908), .A1(n165), .B0(n1480), .B1(n3854), .Y(n2514) );
  OAI22XL U3296 ( .A0(n3905), .A1(n165), .B0(n1481), .B1(n3854), .Y(n2515) );
  OAI22XL U3297 ( .A0(n3920), .A1(n3847), .B0(n1508), .B1(n3848), .Y(n2542) );
  OAI22XL U3298 ( .A0(n3917), .A1(n3847), .B0(n1509), .B1(n3848), .Y(n2543) );
  OAI22XL U3299 ( .A0(n3914), .A1(n3847), .B0(n1510), .B1(n3848), .Y(n2544) );
  OAI22XL U3300 ( .A0(n3911), .A1(n3847), .B0(n1511), .B1(n3848), .Y(n2545) );
  OAI22XL U3301 ( .A0(n3908), .A1(n3846), .B0(n1512), .B1(n3848), .Y(n2546) );
  OAI22XL U3302 ( .A0(n3905), .A1(n3847), .B0(n1513), .B1(n3848), .Y(n2547) );
  OAI22XL U3303 ( .A0(n3921), .A1(n3821), .B0(n1540), .B1(n3822), .Y(n2574) );
  OAI22XL U3304 ( .A0(n3918), .A1(n3821), .B0(n1541), .B1(n3822), .Y(n2575) );
  OAI22XL U3305 ( .A0(n3915), .A1(n3821), .B0(n1542), .B1(n3822), .Y(n2576) );
  OAI22XL U3306 ( .A0(n3912), .A1(n3821), .B0(n1543), .B1(n3822), .Y(n2577) );
  OAI22XL U3307 ( .A0(n3909), .A1(n201), .B0(n1544), .B1(n3822), .Y(n2578) );
  OAI22XL U3308 ( .A0(n3906), .A1(n201), .B0(n1545), .B1(n3822), .Y(n2579) );
  AND4X1 U3309 ( .A(n349), .B(n350), .C(n351), .D(n352), .Y(n129) );
  AOI222XL U3310 ( .A0(dataout[25]), .A1(n252), .B0(N953), .B1(n3775), .C0(
        n3997), .C1(n4011), .Y(n349) );
  AOI222XL U3311 ( .A0(N921), .A1(n253), .B0(N889), .B1(n3778), .C0(N810), 
        .C1(n249), .Y(n350) );
  AOI222XL U3312 ( .A0(N682), .A1(n247), .B0(n2650), .B1(n353), .C0(N228), 
        .C1(n354), .Y(n352) );
  AND4X1 U3313 ( .A(n355), .B(n356), .C(n357), .D(n358), .Y(n130) );
  AOI222XL U3314 ( .A0(dataout[24]), .A1(n3771), .B0(N952), .B1(n3776), .C0(
        n3997), .C1(n2699), .Y(n355) );
  AOI222XL U3315 ( .A0(N920), .A1(n3777), .B0(N888), .B1(n251), .C0(N809), 
        .C1(n3782), .Y(n356) );
  AOI222XL U3316 ( .A0(N681), .A1(n3781), .B0(N197), .B1(n359), .C0(N229), 
        .C1(n360), .Y(n358) );
  AND4X1 U3317 ( .A(n361), .B(n362), .C(n363), .D(n364), .Y(n131) );
  AOI222XL U3318 ( .A0(dataout[23]), .A1(n3772), .B0(N951), .B1(n3776), .C0(
        n3997), .C1(n2725), .Y(n361) );
  AOI222XL U3319 ( .A0(N919), .A1(n253), .B0(N887), .B1(n3778), .C0(N808), 
        .C1(n249), .Y(n362) );
  AOI222XL U3320 ( .A0(N680), .A1(n247), .B0(N198), .B1(n365), .C0(N230), .C1(
        n366), .Y(n364) );
  AND4X1 U3321 ( .A(n367), .B(n368), .C(n369), .D(n370), .Y(n132) );
  AOI222XL U3322 ( .A0(dataout[22]), .A1(n252), .B0(N950), .B1(n3775), .C0(
        n3997), .C1(n2707), .Y(n367) );
  AOI222XL U3323 ( .A0(N918), .A1(n3777), .B0(N886), .B1(n251), .C0(N807), 
        .C1(n3782), .Y(n368) );
  AOI222XL U3324 ( .A0(N679), .A1(n3781), .B0(N199), .B1(n371), .C0(N231), 
        .C1(n372), .Y(n370) );
  AOI222XL U3325 ( .A0(dataout[21]), .A1(n3771), .B0(N949), .B1(n3776), .C0(
        n3997), .C1(n2728), .Y(n373) );
  AOI222XL U3326 ( .A0(N917), .A1(n253), .B0(N885), .B1(n3778), .C0(N806), 
        .C1(n249), .Y(n374) );
  AOI222XL U3327 ( .A0(N678), .A1(n247), .B0(N200), .B1(n377), .C0(N232), .C1(
        n378), .Y(n376) );
  AOI222XL U3328 ( .A0(dataout[20]), .A1(n3772), .B0(N948), .B1(n254), .C0(
        n3997), .C1(n4012), .Y(n379) );
  AOI222XL U3329 ( .A0(N916), .A1(n3777), .B0(N884), .B1(n251), .C0(N805), 
        .C1(n3782), .Y(n380) );
  AOI222XL U3330 ( .A0(N677), .A1(n3781), .B0(n2648), .B1(n383), .C0(N233), 
        .C1(n384), .Y(n382) );
  NOR2X1 U3331 ( .A(\R[3][31] ), .B(n3191), .Y(n3017) );
  NOR2X1 U3332 ( .A(\R[3][30] ), .B(n3191), .Y(n3022) );
  NOR2X1 U3333 ( .A(\R[3][29] ), .B(n3191), .Y(n3027) );
  NOR2X1 U3334 ( .A(\R[3][28] ), .B(n3192), .Y(n3032) );
  NOR2X1 U3335 ( .A(\R[3][27] ), .B(n3192), .Y(n3037) );
  NOR2X1 U3336 ( .A(\R[3][26] ), .B(n3192), .Y(n3042) );
  NOR2X1 U3337 ( .A(\R[3][25] ), .B(n3192), .Y(n3047) );
  NOR2X1 U3338 ( .A(\R[3][24] ), .B(n3193), .Y(n3052) );
  NOR2X1 U3339 ( .A(\R[3][23] ), .B(n3193), .Y(n3057) );
  NOR2X1 U3340 ( .A(\R[3][22] ), .B(n3193), .Y(n3062) );
  NOR2X1 U3341 ( .A(\R[3][21] ), .B(n3193), .Y(n3067) );
  NOR2X1 U3342 ( .A(\R[3][20] ), .B(n3194), .Y(n3072) );
  NOR2X1 U3343 ( .A(\R[3][19] ), .B(n3194), .Y(n3077) );
  NOR2X1 U3344 ( .A(\R[3][18] ), .B(n3194), .Y(n3082) );
  NOR2X1 U3345 ( .A(\R[3][17] ), .B(n3194), .Y(n3087) );
  NOR2X1 U3346 ( .A(\R[3][16] ), .B(n3195), .Y(n3092) );
  NOR2X1 U3347 ( .A(\R[3][15] ), .B(n3195), .Y(n3097) );
  NOR2X1 U3348 ( .A(\R[3][14] ), .B(n3195), .Y(n3102) );
  NOR2X1 U3349 ( .A(\R[3][13] ), .B(n3195), .Y(n3107) );
  NOR2X1 U3350 ( .A(\R[3][12] ), .B(n3196), .Y(n3112) );
  NOR2X1 U3351 ( .A(\R[3][11] ), .B(n3196), .Y(n3117) );
  NOR2X1 U3352 ( .A(\R[3][10] ), .B(n3196), .Y(n3122) );
  NOR2X1 U3353 ( .A(\R[3][9] ), .B(n3196), .Y(n3127) );
  NOR2X1 U3354 ( .A(\R[3][8] ), .B(n3197), .Y(n3132) );
  NOR2X1 U3355 ( .A(\R[3][7] ), .B(n3198), .Y(n3137) );
  NOR2X1 U3356 ( .A(n3212), .B(\R[1][9] ), .Y(n3129) );
  NOR2X1 U3357 ( .A(n3212), .B(\R[1][8] ), .Y(n3134) );
  NOR2X1 U3358 ( .A(n3212), .B(\R[1][7] ), .Y(n3139) );
  AND4X1 U3359 ( .A(instruction[29]), .B(n525), .C(n4001), .D(n3994), .Y(n539)
         );
  AND2X2 U3360 ( .A(n552), .B(instruction[30]), .Y(n543) );
  CLKBUFX3 U3361 ( .A(N47), .Y(n3214) );
  MXI4X1 U3362 ( .A(\R[20][31] ), .B(\R[21][31] ), .C(\R[22][31] ), .D(
        \R[23][31] ), .S0(n3179), .S1(n3209), .Y(n3011) );
  MXI4X1 U3363 ( .A(\R[4][31] ), .B(\R[5][31] ), .C(\R[6][31] ), .D(\R[7][31] ), .S0(n3181), .S1(n3206), .Y(n3015) );
  MXI4X1 U3364 ( .A(\R[20][30] ), .B(\R[21][30] ), .C(\R[22][30] ), .D(
        \R[23][30] ), .S0(n3179), .S1(n3209), .Y(n3003) );
  MXI4X1 U3365 ( .A(\R[4][30] ), .B(\R[5][30] ), .C(\R[6][30] ), .D(\R[7][30] ), .S0(n3179), .S1(n3209), .Y(n3007) );
  MXI4X1 U3366 ( .A(\R[20][29] ), .B(\R[21][29] ), .C(\R[22][29] ), .D(
        \R[23][29] ), .S0(n3179), .S1(n3209), .Y(n2995) );
  MXI4X1 U3367 ( .A(\R[4][29] ), .B(\R[5][29] ), .C(\R[6][29] ), .D(\R[7][29] ), .S0(n3179), .S1(n3209), .Y(n2999) );
  MXI4X1 U3368 ( .A(\R[20][28] ), .B(\R[21][28] ), .C(\R[22][28] ), .D(
        \R[23][28] ), .S0(n3178), .S1(n3209), .Y(n2987) );
  MXI4X1 U3369 ( .A(\R[4][28] ), .B(\R[5][28] ), .C(\R[6][28] ), .D(\R[7][28] ), .S0(n3178), .S1(n3209), .Y(n2991) );
  MXI4X1 U3370 ( .A(\R[20][27] ), .B(\R[21][27] ), .C(\R[22][27] ), .D(
        \R[23][27] ), .S0(n3178), .S1(n3209), .Y(n2979) );
  MXI4X1 U3371 ( .A(\R[4][27] ), .B(\R[5][27] ), .C(\R[6][27] ), .D(\R[7][27] ), .S0(n3178), .S1(n3209), .Y(n2983) );
  MXI4X1 U3372 ( .A(\R[20][26] ), .B(\R[21][26] ), .C(\R[22][26] ), .D(
        \R[23][26] ), .S0(n3178), .S1(n3209), .Y(n2971) );
  MXI4X1 U3373 ( .A(\R[4][26] ), .B(\R[5][26] ), .C(\R[6][26] ), .D(\R[7][26] ), .S0(n3178), .S1(n3209), .Y(n2975) );
  MXI4X1 U3374 ( .A(\R[20][25] ), .B(\R[21][25] ), .C(\R[22][25] ), .D(
        \R[23][25] ), .S0(n3178), .S1(n3209), .Y(n2963) );
  MXI4X1 U3375 ( .A(\R[4][25] ), .B(\R[5][25] ), .C(\R[6][25] ), .D(\R[7][25] ), .S0(n3178), .S1(n3209), .Y(n2967) );
  MXI4X1 U3376 ( .A(\R[20][24] ), .B(\R[21][24] ), .C(\R[22][24] ), .D(
        \R[23][24] ), .S0(n3178), .S1(n3209), .Y(n2955) );
  MXI4X1 U3377 ( .A(\R[4][24] ), .B(\R[5][24] ), .C(\R[6][24] ), .D(\R[7][24] ), .S0(n3178), .S1(n3209), .Y(n2959) );
  MXI4X1 U3378 ( .A(\R[20][23] ), .B(\R[21][23] ), .C(\R[22][23] ), .D(
        \R[23][23] ), .S0(n3178), .S1(n3209), .Y(n2947) );
  MXI4X1 U3379 ( .A(\R[4][23] ), .B(\R[5][23] ), .C(\R[6][23] ), .D(\R[7][23] ), .S0(n3178), .S1(n3209), .Y(n2951) );
  MXI4X1 U3380 ( .A(\R[20][22] ), .B(\R[21][22] ), .C(\R[22][22] ), .D(
        \R[23][22] ), .S0(n3178), .S1(n3208), .Y(n2939) );
  MXI4X1 U3381 ( .A(\R[4][22] ), .B(\R[5][22] ), .C(\R[6][22] ), .D(\R[7][22] ), .S0(n3178), .S1(n3209), .Y(n2943) );
  MXI4X1 U3382 ( .A(\R[20][21] ), .B(\R[21][21] ), .C(\R[22][21] ), .D(
        \R[23][21] ), .S0(n3178), .S1(n3208), .Y(n2931) );
  MXI4X1 U3383 ( .A(\R[4][21] ), .B(\R[5][21] ), .C(\R[6][21] ), .D(\R[7][21] ), .S0(n3178), .S1(n3208), .Y(n2935) );
  MXI4X1 U3384 ( .A(\R[20][15] ), .B(\R[21][15] ), .C(\R[22][15] ), .D(
        \R[23][15] ), .S0(n3181), .S1(n3208), .Y(n2883) );
  MXI4X1 U3385 ( .A(\R[4][15] ), .B(\R[5][15] ), .C(\R[6][15] ), .D(\R[7][15] ), .S0(n3180), .S1(n3208), .Y(n2887) );
  MXI4X1 U3386 ( .A(\R[20][14] ), .B(\R[21][14] ), .C(\R[22][14] ), .D(
        \R[23][14] ), .S0(n3181), .S1(n3208), .Y(n2875) );
  MXI4X1 U3387 ( .A(\R[4][14] ), .B(\R[5][14] ), .C(\R[6][14] ), .D(\R[7][14] ), .S0(n3181), .S1(n3208), .Y(n2879) );
  MXI4X1 U3388 ( .A(\R[20][13] ), .B(\R[21][13] ), .C(\R[22][13] ), .D(
        \R[23][13] ), .S0(n3180), .S1(n3208), .Y(n2867) );
  MXI4X1 U3389 ( .A(\R[4][13] ), .B(\R[5][13] ), .C(\R[6][13] ), .D(\R[7][13] ), .S0(n3181), .S1(n3208), .Y(n2871) );
  MXI4X1 U3390 ( .A(\R[20][11] ), .B(\R[21][11] ), .C(\R[22][11] ), .D(
        \R[23][11] ), .S0(n3180), .S1(n3207), .Y(n2851) );
  MXI4X1 U3391 ( .A(\R[4][11] ), .B(\R[5][11] ), .C(\R[6][11] ), .D(\R[7][11] ), .S0(n3180), .S1(n3207), .Y(n2855) );
  MXI4X1 U3392 ( .A(\R[20][10] ), .B(\R[21][10] ), .C(\R[22][10] ), .D(
        \R[23][10] ), .S0(n3180), .S1(n3207), .Y(n2843) );
  MXI4X1 U3393 ( .A(\R[4][10] ), .B(\R[5][10] ), .C(\R[6][10] ), .D(\R[7][10] ), .S0(n3180), .S1(n3207), .Y(n2847) );
  MXI4X1 U3394 ( .A(\R[20][9] ), .B(\R[21][9] ), .C(\R[22][9] ), .D(\R[23][9] ), .S0(n3180), .S1(n3207), .Y(n2835) );
  MXI4X1 U3395 ( .A(\R[4][9] ), .B(\R[5][9] ), .C(\R[6][9] ), .D(\R[7][9] ), 
        .S0(n3180), .S1(n3207), .Y(n2839) );
  MXI4X1 U3396 ( .A(\R[20][8] ), .B(\R[21][8] ), .C(\R[22][8] ), .D(\R[23][8] ), .S0(n3180), .S1(n3207), .Y(n2827) );
  MXI4X1 U3397 ( .A(\R[4][8] ), .B(\R[5][8] ), .C(\R[6][8] ), .D(\R[7][8] ), 
        .S0(n3180), .S1(n3207), .Y(n2831) );
  MXI4X1 U3398 ( .A(\R[20][7] ), .B(\R[21][7] ), .C(\R[22][7] ), .D(\R[23][7] ), .S0(n3180), .S1(n3207), .Y(n2819) );
  MXI4X1 U3399 ( .A(\R[4][7] ), .B(\R[5][7] ), .C(\R[6][7] ), .D(\R[7][7] ), 
        .S0(n3180), .S1(n3207), .Y(n2823) );
  MXI4X1 U3400 ( .A(\R[20][20] ), .B(\R[21][20] ), .C(\R[22][20] ), .D(
        \R[23][20] ), .S0(n3177), .S1(n3208), .Y(n2923) );
  MXI4X1 U3401 ( .A(\R[4][20] ), .B(\R[5][20] ), .C(\R[6][20] ), .D(\R[7][20] ), .S0(n3177), .S1(n3208), .Y(n2927) );
  MXI4X1 U3402 ( .A(\R[20][19] ), .B(\R[21][19] ), .C(\R[22][19] ), .D(
        \R[23][19] ), .S0(n3177), .S1(n3208), .Y(n2915) );
  MXI4X1 U3403 ( .A(\R[4][19] ), .B(\R[5][19] ), .C(\R[6][19] ), .D(\R[7][19] ), .S0(n3177), .S1(n3208), .Y(n2919) );
  MXI4X1 U3404 ( .A(\R[20][18] ), .B(\R[21][18] ), .C(\R[22][18] ), .D(
        \R[23][18] ), .S0(n3177), .S1(n3208), .Y(n2907) );
  MXI4X1 U3405 ( .A(\R[4][18] ), .B(\R[5][18] ), .C(\R[6][18] ), .D(\R[7][18] ), .S0(n3177), .S1(n3208), .Y(n2911) );
  MXI4X1 U3406 ( .A(\R[20][17] ), .B(\R[21][17] ), .C(\R[22][17] ), .D(
        \R[23][17] ), .S0(n3177), .S1(n3208), .Y(n2899) );
  MXI4X1 U3407 ( .A(\R[4][17] ), .B(\R[5][17] ), .C(\R[6][17] ), .D(\R[7][17] ), .S0(n3177), .S1(n3208), .Y(n2903) );
  MXI4X1 U3408 ( .A(\R[20][16] ), .B(\R[21][16] ), .C(\R[22][16] ), .D(
        \R[23][16] ), .S0(n3177), .S1(n3208), .Y(n2891) );
  MXI4X1 U3409 ( .A(\R[4][16] ), .B(\R[5][16] ), .C(\R[6][16] ), .D(\R[7][16] ), .S0(n3177), .S1(n3208), .Y(n2895) );
  MXI4X1 U3410 ( .A(\R[16][31] ), .B(\R[17][31] ), .C(\R[18][31] ), .D(
        \R[19][31] ), .S0(n3179), .S1(n3209), .Y(n3009) );
  MXI4X1 U3411 ( .A(\R[16][30] ), .B(\R[17][30] ), .C(\R[18][30] ), .D(
        \R[19][30] ), .S0(n3179), .S1(n3209), .Y(n3001) );
  MXI4X1 U3412 ( .A(\R[16][29] ), .B(\R[17][29] ), .C(\R[18][29] ), .D(
        \R[19][29] ), .S0(n3179), .S1(n3209), .Y(n2993) );
  MXI4X1 U3413 ( .A(\R[16][28] ), .B(\R[17][28] ), .C(\R[18][28] ), .D(
        \R[19][28] ), .S0(n3178), .S1(n3209), .Y(n2985) );
  MXI4X1 U3414 ( .A(\R[16][27] ), .B(\R[17][27] ), .C(\R[18][27] ), .D(
        \R[19][27] ), .S0(n3178), .S1(n3209), .Y(n2977) );
  MXI4X1 U3415 ( .A(\R[16][26] ), .B(\R[17][26] ), .C(\R[18][26] ), .D(
        \R[19][26] ), .S0(n3178), .S1(n3209), .Y(n2969) );
  MXI4X1 U3416 ( .A(\R[16][25] ), .B(\R[17][25] ), .C(\R[18][25] ), .D(
        \R[19][25] ), .S0(n3178), .S1(n3209), .Y(n2961) );
  MXI4X1 U3417 ( .A(\R[16][24] ), .B(\R[17][24] ), .C(\R[18][24] ), .D(
        \R[19][24] ), .S0(n3178), .S1(n3209), .Y(n2953) );
  MXI4X1 U3418 ( .A(\R[16][23] ), .B(\R[17][23] ), .C(\R[18][23] ), .D(
        \R[19][23] ), .S0(n3178), .S1(n3209), .Y(n2945) );
  MXI4X1 U3419 ( .A(\R[16][22] ), .B(\R[17][22] ), .C(\R[18][22] ), .D(
        \R[19][22] ), .S0(n3178), .S1(n3208), .Y(n2937) );
  MXI4X1 U3420 ( .A(\R[16][21] ), .B(\R[17][21] ), .C(\R[18][21] ), .D(
        \R[19][21] ), .S0(n3178), .S1(n3208), .Y(n2929) );
  MXI4X1 U3421 ( .A(\R[16][15] ), .B(\R[17][15] ), .C(\R[18][15] ), .D(
        \R[19][15] ), .S0(n3181), .S1(n3208), .Y(n2881) );
  MXI4X1 U3422 ( .A(\R[16][14] ), .B(\R[17][14] ), .C(\R[18][14] ), .D(
        \R[19][14] ), .S0(n3181), .S1(n3208), .Y(n2873) );
  MXI4X1 U3423 ( .A(\R[16][13] ), .B(\R[17][13] ), .C(\R[18][13] ), .D(
        \R[19][13] ), .S0(n3180), .S1(n3208), .Y(n2865) );
  MXI4X1 U3424 ( .A(\R[16][12] ), .B(\R[17][12] ), .C(\R[18][12] ), .D(
        \R[19][12] ), .S0(n3180), .S1(n3207), .Y(n2857) );
  MXI4X1 U3425 ( .A(\R[16][11] ), .B(\R[17][11] ), .C(\R[18][11] ), .D(
        \R[19][11] ), .S0(n3180), .S1(n3207), .Y(n2849) );
  MXI4X1 U3426 ( .A(\R[16][10] ), .B(\R[17][10] ), .C(\R[18][10] ), .D(
        \R[19][10] ), .S0(n3180), .S1(n3207), .Y(n2841) );
  MXI4X1 U3427 ( .A(\R[16][9] ), .B(\R[17][9] ), .C(\R[18][9] ), .D(\R[19][9] ), .S0(n3180), .S1(n3207), .Y(n2833) );
  MXI4X1 U3428 ( .A(\R[16][8] ), .B(\R[17][8] ), .C(\R[18][8] ), .D(\R[19][8] ), .S0(n3180), .S1(n3207), .Y(n2825) );
  MXI4X1 U3429 ( .A(\R[16][7] ), .B(\R[17][7] ), .C(\R[18][7] ), .D(\R[19][7] ), .S0(n3180), .S1(n3207), .Y(n2817) );
  MXI4X1 U3430 ( .A(\R[16][20] ), .B(\R[17][20] ), .C(\R[18][20] ), .D(
        \R[19][20] ), .S0(n3177), .S1(n3208), .Y(n2921) );
  MXI4X1 U3431 ( .A(\R[16][19] ), .B(\R[17][19] ), .C(\R[18][19] ), .D(
        \R[19][19] ), .S0(n3177), .S1(n3208), .Y(n2913) );
  MXI4X1 U3432 ( .A(\R[16][18] ), .B(\R[17][18] ), .C(\R[18][18] ), .D(
        \R[19][18] ), .S0(n3177), .S1(n3208), .Y(n2905) );
  MXI4X1 U3433 ( .A(\R[16][17] ), .B(\R[17][17] ), .C(\R[18][17] ), .D(
        \R[19][17] ), .S0(n3177), .S1(n3208), .Y(n2897) );
  MXI4X1 U3434 ( .A(\R[16][16] ), .B(\R[17][16] ), .C(\R[18][16] ), .D(
        \R[19][16] ), .S0(n3177), .S1(n3208), .Y(n2889) );
  MXI4X1 U3435 ( .A(\R[24][31] ), .B(\R[25][31] ), .C(\R[26][31] ), .D(
        \R[27][31] ), .S0(n3179), .S1(n3209), .Y(n3010) );
  MXI4X1 U3436 ( .A(\R[8][31] ), .B(\R[9][31] ), .C(\R[10][31] ), .D(
        \R[11][31] ), .S0(n3178), .S1(n3209), .Y(n3014) );
  MXI4X1 U3437 ( .A(\R[24][30] ), .B(\R[25][30] ), .C(\R[26][30] ), .D(
        \R[27][30] ), .S0(n3179), .S1(n3209), .Y(n3002) );
  MXI4X1 U3438 ( .A(\R[8][30] ), .B(\R[9][30] ), .C(\R[10][30] ), .D(
        \R[11][30] ), .S0(n3179), .S1(n3209), .Y(n3006) );
  MXI4X1 U3439 ( .A(\R[24][29] ), .B(\R[25][29] ), .C(\R[26][29] ), .D(
        \R[27][29] ), .S0(n3179), .S1(n3209), .Y(n2994) );
  MXI4X1 U3440 ( .A(\R[8][29] ), .B(\R[9][29] ), .C(\R[10][29] ), .D(
        \R[11][29] ), .S0(n3179), .S1(n3209), .Y(n2998) );
  MXI4X1 U3441 ( .A(\R[24][28] ), .B(\R[25][28] ), .C(\R[26][28] ), .D(
        \R[27][28] ), .S0(n3178), .S1(n3209), .Y(n2986) );
  MXI4X1 U3442 ( .A(\R[8][28] ), .B(\R[9][28] ), .C(\R[10][28] ), .D(
        \R[11][28] ), .S0(n3178), .S1(n3209), .Y(n2990) );
  MXI4X1 U3443 ( .A(\R[24][27] ), .B(\R[25][27] ), .C(\R[26][27] ), .D(
        \R[27][27] ), .S0(n3178), .S1(n3209), .Y(n2978) );
  MXI4X1 U3444 ( .A(\R[8][27] ), .B(\R[9][27] ), .C(\R[10][27] ), .D(
        \R[11][27] ), .S0(n3178), .S1(n3209), .Y(n2982) );
  MXI4X1 U3445 ( .A(\R[24][26] ), .B(\R[25][26] ), .C(\R[26][26] ), .D(
        \R[27][26] ), .S0(n3178), .S1(n3209), .Y(n2970) );
  MXI4X1 U3446 ( .A(\R[8][26] ), .B(\R[9][26] ), .C(\R[10][26] ), .D(
        \R[11][26] ), .S0(n3178), .S1(n3209), .Y(n2974) );
  MXI4X1 U3447 ( .A(\R[24][25] ), .B(\R[25][25] ), .C(\R[26][25] ), .D(
        \R[27][25] ), .S0(n3178), .S1(n3209), .Y(n2962) );
  MXI4X1 U3448 ( .A(\R[8][25] ), .B(\R[9][25] ), .C(\R[10][25] ), .D(
        \R[11][25] ), .S0(n3178), .S1(n3209), .Y(n2966) );
  MXI4X1 U3449 ( .A(\R[24][24] ), .B(\R[25][24] ), .C(\R[26][24] ), .D(
        \R[27][24] ), .S0(n3178), .S1(n3209), .Y(n2954) );
  MXI4X1 U3450 ( .A(\R[8][24] ), .B(\R[9][24] ), .C(\R[10][24] ), .D(
        \R[11][24] ), .S0(n3178), .S1(n3209), .Y(n2958) );
  MXI4X1 U3451 ( .A(\R[24][23] ), .B(\R[25][23] ), .C(\R[26][23] ), .D(
        \R[27][23] ), .S0(n3178), .S1(n3209), .Y(n2946) );
  MXI4X1 U3452 ( .A(\R[8][23] ), .B(\R[9][23] ), .C(\R[10][23] ), .D(
        \R[11][23] ), .S0(n3178), .S1(n3209), .Y(n2950) );
  MXI4X1 U3453 ( .A(\R[24][22] ), .B(\R[25][22] ), .C(\R[26][22] ), .D(
        \R[27][22] ), .S0(n3178), .S1(n3208), .Y(n2938) );
  MXI4X1 U3454 ( .A(\R[8][22] ), .B(\R[9][22] ), .C(\R[10][22] ), .D(
        \R[11][22] ), .S0(n3178), .S1(n3209), .Y(n2942) );
  MXI4X1 U3455 ( .A(\R[24][21] ), .B(\R[25][21] ), .C(\R[26][21] ), .D(
        \R[27][21] ), .S0(n3178), .S1(n3208), .Y(n2930) );
  MXI4X1 U3456 ( .A(\R[8][21] ), .B(\R[9][21] ), .C(\R[10][21] ), .D(
        \R[11][21] ), .S0(n3178), .S1(n3208), .Y(n2934) );
  MXI4X1 U3457 ( .A(\R[24][15] ), .B(\R[25][15] ), .C(\R[26][15] ), .D(
        \R[27][15] ), .S0(n3181), .S1(n3208), .Y(n2882) );
  MXI4X1 U3458 ( .A(\R[8][15] ), .B(\R[9][15] ), .C(\R[10][15] ), .D(
        \R[11][15] ), .S0(n3181), .S1(n3208), .Y(n2886) );
  MXI4X1 U3459 ( .A(\R[24][14] ), .B(\R[25][14] ), .C(\R[26][14] ), .D(
        \R[27][14] ), .S0(n3181), .S1(n3208), .Y(n2874) );
  MXI4X1 U3460 ( .A(\R[8][14] ), .B(\R[9][14] ), .C(\R[10][14] ), .D(
        \R[11][14] ), .S0(n3181), .S1(n3208), .Y(n2878) );
  MXI4X1 U3461 ( .A(\R[24][13] ), .B(\R[25][13] ), .C(\R[26][13] ), .D(
        \R[27][13] ), .S0(n3180), .S1(n3207), .Y(n2866) );
  MXI4X1 U3462 ( .A(\R[8][13] ), .B(\R[9][13] ), .C(\R[10][13] ), .D(
        \R[11][13] ), .S0(n3180), .S1(n3208), .Y(n2870) );
  MXI4X1 U3463 ( .A(\R[8][10] ), .B(\R[9][10] ), .C(\R[10][10] ), .D(
        \R[11][10] ), .S0(n3180), .S1(n3207), .Y(n2846) );
  MXI4X1 U3464 ( .A(\R[24][9] ), .B(\R[25][9] ), .C(\R[26][9] ), .D(\R[27][9] ), .S0(n3180), .S1(n3207), .Y(n2834) );
  MXI4X1 U3465 ( .A(\R[8][9] ), .B(\R[9][9] ), .C(\R[10][9] ), .D(\R[11][9] ), 
        .S0(n3180), .S1(n3207), .Y(n2838) );
  MXI4X1 U3466 ( .A(\R[24][8] ), .B(\R[25][8] ), .C(\R[26][8] ), .D(\R[27][8] ), .S0(n3180), .S1(n3207), .Y(n2826) );
  MXI4X1 U3467 ( .A(\R[8][8] ), .B(\R[9][8] ), .C(\R[10][8] ), .D(\R[11][8] ), 
        .S0(n3180), .S1(n3207), .Y(n2830) );
  MXI4X1 U3468 ( .A(\R[24][7] ), .B(\R[25][7] ), .C(\R[26][7] ), .D(\R[27][7] ), .S0(n3180), .S1(n3207), .Y(n2818) );
  MXI4X1 U3469 ( .A(\R[8][7] ), .B(\R[9][7] ), .C(\R[10][7] ), .D(\R[11][7] ), 
        .S0(n3180), .S1(n3207), .Y(n2822) );
  MXI4X1 U3470 ( .A(\R[24][20] ), .B(\R[25][20] ), .C(\R[26][20] ), .D(
        \R[27][20] ), .S0(n3177), .S1(n3208), .Y(n2922) );
  MXI4X1 U3471 ( .A(\R[8][20] ), .B(\R[9][20] ), .C(\R[10][20] ), .D(
        \R[11][20] ), .S0(n3177), .S1(n3208), .Y(n2926) );
  MXI4X1 U3472 ( .A(\R[24][19] ), .B(\R[25][19] ), .C(\R[26][19] ), .D(
        \R[27][19] ), .S0(n3177), .S1(n3208), .Y(n2914) );
  MXI4X1 U3473 ( .A(\R[8][19] ), .B(\R[9][19] ), .C(\R[10][19] ), .D(
        \R[11][19] ), .S0(n3177), .S1(n3208), .Y(n2918) );
  MXI4X1 U3474 ( .A(\R[24][18] ), .B(\R[25][18] ), .C(\R[26][18] ), .D(
        \R[27][18] ), .S0(n3177), .S1(n3208), .Y(n2906) );
  MXI4X1 U3475 ( .A(\R[8][18] ), .B(\R[9][18] ), .C(\R[10][18] ), .D(
        \R[11][18] ), .S0(n3177), .S1(n3208), .Y(n2910) );
  MXI4X1 U3476 ( .A(\R[24][17] ), .B(\R[25][17] ), .C(\R[26][17] ), .D(
        \R[27][17] ), .S0(n3177), .S1(n3208), .Y(n2898) );
  MXI4X1 U3477 ( .A(\R[8][17] ), .B(\R[9][17] ), .C(\R[10][17] ), .D(
        \R[11][17] ), .S0(n3177), .S1(n3208), .Y(n2902) );
  MXI4X1 U3478 ( .A(\R[24][16] ), .B(\R[25][16] ), .C(\R[26][16] ), .D(
        \R[27][16] ), .S0(n3177), .S1(n3208), .Y(n2890) );
  MXI4X1 U3479 ( .A(\R[8][16] ), .B(\R[9][16] ), .C(\R[10][16] ), .D(
        \R[11][16] ), .S0(n3177), .S1(n3208), .Y(n2894) );
  MXI4X1 U3480 ( .A(\R[28][31] ), .B(\R[29][31] ), .C(\R[30][31] ), .D(
        \R[31][31] ), .S0(n3179), .S1(n3209), .Y(n3012) );
  MXI4X1 U3481 ( .A(\R[12][31] ), .B(\R[13][31] ), .C(\R[14][31] ), .D(
        \R[15][31] ), .S0(n3179), .S1(n3209), .Y(n3016) );
  MXI4X1 U3482 ( .A(\R[28][30] ), .B(\R[29][30] ), .C(\R[30][30] ), .D(
        \R[31][30] ), .S0(n3179), .S1(n3209), .Y(n3004) );
  MXI4X1 U3483 ( .A(\R[12][30] ), .B(\R[13][30] ), .C(\R[14][30] ), .D(
        \R[15][30] ), .S0(n3179), .S1(n3209), .Y(n3008) );
  MXI4X1 U3484 ( .A(\R[28][29] ), .B(\R[29][29] ), .C(\R[30][29] ), .D(
        \R[31][29] ), .S0(n3178), .S1(n3209), .Y(n2996) );
  MXI4X1 U3485 ( .A(\R[12][29] ), .B(\R[13][29] ), .C(\R[14][29] ), .D(
        \R[15][29] ), .S0(n3179), .S1(n3209), .Y(n3000) );
  MXI4X1 U3486 ( .A(\R[28][28] ), .B(\R[29][28] ), .C(\R[30][28] ), .D(
        \R[31][28] ), .S0(n3178), .S1(n3209), .Y(n2988) );
  MXI4X1 U3487 ( .A(\R[12][28] ), .B(\R[13][28] ), .C(\R[14][28] ), .D(
        \R[15][28] ), .S0(n3178), .S1(n3209), .Y(n2992) );
  MXI4X1 U3488 ( .A(\R[28][27] ), .B(\R[29][27] ), .C(\R[30][27] ), .D(
        \R[31][27] ), .S0(n3178), .S1(n3209), .Y(n2980) );
  MXI4X1 U3489 ( .A(\R[12][27] ), .B(\R[13][27] ), .C(\R[14][27] ), .D(
        \R[15][27] ), .S0(n3178), .S1(n3209), .Y(n2984) );
  MXI4X1 U3490 ( .A(\R[28][26] ), .B(\R[29][26] ), .C(\R[30][26] ), .D(
        \R[31][26] ), .S0(n3178), .S1(n3209), .Y(n2972) );
  MXI4X1 U3491 ( .A(\R[12][26] ), .B(\R[13][26] ), .C(\R[14][26] ), .D(
        \R[15][26] ), .S0(n3178), .S1(n3209), .Y(n2976) );
  MXI4X1 U3492 ( .A(\R[28][25] ), .B(\R[29][25] ), .C(\R[30][25] ), .D(
        \R[31][25] ), .S0(n3178), .S1(n3209), .Y(n2964) );
  MXI4X1 U3493 ( .A(\R[12][25] ), .B(\R[13][25] ), .C(\R[14][25] ), .D(
        \R[15][25] ), .S0(n3178), .S1(n3209), .Y(n2968) );
  MXI4X1 U3494 ( .A(\R[28][24] ), .B(\R[29][24] ), .C(\R[30][24] ), .D(
        \R[31][24] ), .S0(n3178), .S1(n3209), .Y(n2956) );
  MXI4X1 U3495 ( .A(\R[12][24] ), .B(\R[13][24] ), .C(\R[14][24] ), .D(
        \R[15][24] ), .S0(n3178), .S1(n3209), .Y(n2960) );
  MXI4X1 U3496 ( .A(\R[28][23] ), .B(\R[29][23] ), .C(\R[30][23] ), .D(
        \R[31][23] ), .S0(n3178), .S1(n3209), .Y(n2948) );
  MXI4X1 U3497 ( .A(\R[12][23] ), .B(\R[13][23] ), .C(\R[14][23] ), .D(
        \R[15][23] ), .S0(n3178), .S1(n3209), .Y(n2952) );
  MXI4X1 U3498 ( .A(\R[28][22] ), .B(\R[29][22] ), .C(\R[30][22] ), .D(
        \R[31][22] ), .S0(n3178), .S1(n3208), .Y(n2940) );
  MXI4X1 U3499 ( .A(\R[12][22] ), .B(\R[13][22] ), .C(\R[14][22] ), .D(
        \R[15][22] ), .S0(n3178), .S1(n3209), .Y(n2944) );
  MXI4X1 U3500 ( .A(\R[28][21] ), .B(\R[29][21] ), .C(\R[30][21] ), .D(
        \R[31][21] ), .S0(n3178), .S1(n3208), .Y(n2932) );
  MXI4X1 U3501 ( .A(\R[12][21] ), .B(\R[13][21] ), .C(\R[14][21] ), .D(
        \R[15][21] ), .S0(n3178), .S1(n3208), .Y(n2936) );
  MXI4X1 U3502 ( .A(\R[28][15] ), .B(\R[29][15] ), .C(\R[30][15] ), .D(
        \R[31][15] ), .S0(n3181), .S1(n3208), .Y(n2884) );
  MXI4X1 U3503 ( .A(\R[12][15] ), .B(\R[13][15] ), .C(\R[14][15] ), .D(
        \R[15][15] ), .S0(n3181), .S1(n3208), .Y(n2888) );
  MXI4X1 U3504 ( .A(\R[28][14] ), .B(\R[29][14] ), .C(\R[30][14] ), .D(
        \R[31][14] ), .S0(n3181), .S1(n3208), .Y(n2876) );
  MXI4X1 U3505 ( .A(\R[12][14] ), .B(\R[13][14] ), .C(\R[14][14] ), .D(
        \R[15][14] ), .S0(n3181), .S1(n3208), .Y(n2880) );
  MXI4X1 U3506 ( .A(\R[28][13] ), .B(\R[29][13] ), .C(\R[30][13] ), .D(
        \R[31][13] ), .S0(n3180), .S1(n3207), .Y(n2868) );
  MXI4X1 U3507 ( .A(\R[12][13] ), .B(\R[13][13] ), .C(\R[14][13] ), .D(
        \R[15][13] ), .S0(n3180), .S1(n3208), .Y(n2872) );
  MXI4X1 U3508 ( .A(\R[28][12] ), .B(\R[29][12] ), .C(\R[30][12] ), .D(
        \R[31][12] ), .S0(n3180), .S1(n3207), .Y(n2860) );
  MXI4X1 U3509 ( .A(\R[12][12] ), .B(\R[13][12] ), .C(\R[14][12] ), .D(
        \R[15][12] ), .S0(n3180), .S1(n3207), .Y(n2864) );
  MXI4X1 U3510 ( .A(\R[28][11] ), .B(\R[29][11] ), .C(\R[30][11] ), .D(
        \R[31][11] ), .S0(n3180), .S1(n3207), .Y(n2852) );
  MXI4X1 U3511 ( .A(\R[12][11] ), .B(\R[13][11] ), .C(\R[14][11] ), .D(
        \R[15][11] ), .S0(n3180), .S1(n3207), .Y(n2856) );
  MXI4X1 U3512 ( .A(\R[28][10] ), .B(\R[29][10] ), .C(\R[30][10] ), .D(
        \R[31][10] ), .S0(n3180), .S1(n3207), .Y(n2844) );
  MXI4X1 U3513 ( .A(\R[12][10] ), .B(\R[13][10] ), .C(\R[14][10] ), .D(
        \R[15][10] ), .S0(n3180), .S1(n3207), .Y(n2848) );
  MXI4X1 U3514 ( .A(\R[28][9] ), .B(\R[29][9] ), .C(\R[30][9] ), .D(\R[31][9] ), .S0(n3180), .S1(n3207), .Y(n2836) );
  MXI4X1 U3515 ( .A(\R[12][9] ), .B(\R[13][9] ), .C(\R[14][9] ), .D(\R[15][9] ), .S0(n3180), .S1(n3207), .Y(n2840) );
  MXI4X1 U3516 ( .A(\R[28][8] ), .B(\R[29][8] ), .C(\R[30][8] ), .D(\R[31][8] ), .S0(n3180), .S1(n3207), .Y(n2828) );
  MXI4X1 U3517 ( .A(\R[12][8] ), .B(\R[13][8] ), .C(\R[14][8] ), .D(\R[15][8] ), .S0(n3180), .S1(n3207), .Y(n2832) );
  MXI4X1 U3518 ( .A(\R[28][7] ), .B(\R[29][7] ), .C(\R[30][7] ), .D(\R[31][7] ), .S0(n3180), .S1(n3207), .Y(n2820) );
  MXI4X1 U3519 ( .A(\R[12][7] ), .B(\R[13][7] ), .C(\R[14][7] ), .D(\R[15][7] ), .S0(n3180), .S1(n3207), .Y(n2824) );
  MXI4X1 U3520 ( .A(\R[28][20] ), .B(\R[29][20] ), .C(\R[30][20] ), .D(
        \R[31][20] ), .S0(n3177), .S1(n3208), .Y(n2924) );
  MXI4X1 U3521 ( .A(\R[12][20] ), .B(\R[13][20] ), .C(\R[14][20] ), .D(
        \R[15][20] ), .S0(n3177), .S1(n3208), .Y(n2928) );
  MXI4X1 U3522 ( .A(\R[28][19] ), .B(\R[29][19] ), .C(\R[30][19] ), .D(
        \R[31][19] ), .S0(n3177), .S1(n3208), .Y(n2916) );
  MXI4X1 U3523 ( .A(\R[12][19] ), .B(\R[13][19] ), .C(\R[14][19] ), .D(
        \R[15][19] ), .S0(n3177), .S1(n3208), .Y(n2920) );
  MXI4X1 U3524 ( .A(\R[28][18] ), .B(\R[29][18] ), .C(\R[30][18] ), .D(
        \R[31][18] ), .S0(n3177), .S1(n3208), .Y(n2908) );
  MXI4X1 U3525 ( .A(\R[12][18] ), .B(\R[13][18] ), .C(\R[14][18] ), .D(
        \R[15][18] ), .S0(n3177), .S1(n3208), .Y(n2912) );
  MXI4X1 U3526 ( .A(\R[28][17] ), .B(\R[29][17] ), .C(\R[30][17] ), .D(
        \R[31][17] ), .S0(n3177), .S1(n3208), .Y(n2900) );
  MXI4X1 U3527 ( .A(\R[12][17] ), .B(\R[13][17] ), .C(\R[14][17] ), .D(
        \R[15][17] ), .S0(n3177), .S1(n3208), .Y(n2904) );
  MXI4X1 U3528 ( .A(\R[28][16] ), .B(\R[29][16] ), .C(\R[30][16] ), .D(
        \R[31][16] ), .S0(n3177), .S1(n3208), .Y(n2892) );
  MXI4X1 U3529 ( .A(\R[12][16] ), .B(\R[13][16] ), .C(\R[14][16] ), .D(
        \R[15][16] ), .S0(n3177), .S1(n3208), .Y(n2896) );
  CLKBUFX3 U3530 ( .A(N46), .Y(n3185) );
  CLKBUFX3 U3531 ( .A(N49), .Y(n3230) );
  CLKBUFX3 U3532 ( .A(N49), .Y(n3229) );
  OAI221XL U3533 ( .A0(n2738), .A1(n3783), .B0(n1566), .B1(n4045), .C0(n491), 
        .Y(n2600) );
  AOI22X1 U3534 ( .A0(N283), .A1(n3789), .B0(N1022), .B1(n3785), .Y(n491) );
  OAI221XL U3535 ( .A0(n2696), .A1(n478), .B0(n1567), .B1(n4045), .C0(n492), 
        .Y(n2601) );
  OAI221XL U3536 ( .A0(n4009), .A1(n3783), .B0(n1596), .B1(n4045), .C0(n489), 
        .Y(n2630) );
  OAI221XL U3537 ( .A0(n2735), .A1(n478), .B0(n1607), .B1(n4045), .C0(n488), 
        .Y(n2631) );
  AOI22X1 U3538 ( .A0(N285), .A1(n3789), .B0(N1024), .B1(n3786), .Y(n488) );
  NAND2X1 U3539 ( .A(n3056), .B(n3055), .Y(n2957) );
  NOR2X1 U3540 ( .A(n3054), .B(n3053), .Y(n3056) );
  MXI2X1 U3541 ( .A(n1509), .B(n3052), .S0(n3182), .Y(n3055) );
  NOR2X1 U3542 ( .A(n3210), .B(\R[1][24] ), .Y(n3054) );
  NAND2X1 U3543 ( .A(n3066), .B(n3065), .Y(n2941) );
  NOR2X1 U3544 ( .A(n3064), .B(n3063), .Y(n3066) );
  MXI2X1 U3545 ( .A(n1511), .B(n3062), .S0(n3182), .Y(n3065) );
  NOR2X1 U3546 ( .A(n3210), .B(\R[1][22] ), .Y(n3064) );
  NAND2X1 U3547 ( .A(n3071), .B(n3070), .Y(n2933) );
  NOR2X1 U3548 ( .A(n3069), .B(n3068), .Y(n3071) );
  MXI2X1 U3549 ( .A(n1512), .B(n3067), .S0(n3182), .Y(n3070) );
  NOR2X1 U3550 ( .A(n3210), .B(\R[1][21] ), .Y(n3069) );
  NAND2X1 U3551 ( .A(n3076), .B(n3075), .Y(n2925) );
  NOR2X1 U3552 ( .A(n3074), .B(n3073), .Y(n3076) );
  MXI2X1 U3553 ( .A(n1513), .B(n3072), .S0(n3182), .Y(n3075) );
  NOR2X1 U3554 ( .A(n3210), .B(\R[1][20] ), .Y(n3074) );
  NAND2X1 U3555 ( .A(n3081), .B(n3080), .Y(n2917) );
  NOR2X1 U3556 ( .A(n3079), .B(n3078), .Y(n3081) );
  MXI2X1 U3557 ( .A(n1514), .B(n3077), .S0(n3182), .Y(n3080) );
  NOR2X1 U3558 ( .A(n3211), .B(\R[1][19] ), .Y(n3079) );
  NAND2X1 U3559 ( .A(n3086), .B(n3085), .Y(n2909) );
  NOR2X1 U3560 ( .A(n3084), .B(n3083), .Y(n3086) );
  MXI2X1 U3561 ( .A(n1515), .B(n3082), .S0(n3182), .Y(n3085) );
  NOR2X1 U3562 ( .A(n3211), .B(\R[1][18] ), .Y(n3084) );
  NAND2X1 U3563 ( .A(n3096), .B(n3095), .Y(n2893) );
  NOR2X1 U3564 ( .A(n3094), .B(n3093), .Y(n3096) );
  MXI2X1 U3565 ( .A(n1517), .B(n3092), .S0(n3182), .Y(n3095) );
  NOR2X1 U3566 ( .A(n3211), .B(\R[1][16] ), .Y(n3094) );
  NAND2X1 U3567 ( .A(n3101), .B(n3100), .Y(n2885) );
  NOR2X1 U3568 ( .A(n3099), .B(n3098), .Y(n3101) );
  MXI2X1 U3569 ( .A(n1518), .B(n3097), .S0(n3182), .Y(n3100) );
  NOR2X1 U3570 ( .A(n3211), .B(\R[1][15] ), .Y(n3099) );
  NAND2X1 U3571 ( .A(n3021), .B(n3020), .Y(n3013) );
  NOR2X1 U3572 ( .A(n3019), .B(n3018), .Y(n3021) );
  MXI2X1 U3573 ( .A(n1502), .B(n3017), .S0(n3184), .Y(n3020) );
  NOR2X1 U3574 ( .A(n3213), .B(\R[1][31] ), .Y(n3019) );
  NAND2X1 U3575 ( .A(n3026), .B(n3025), .Y(n3005) );
  NOR2X1 U3576 ( .A(n3024), .B(n3023), .Y(n3026) );
  MXI2X1 U3577 ( .A(n1503), .B(n3022), .S0(n3184), .Y(n3025) );
  NOR2X1 U3578 ( .A(n3206), .B(\R[1][30] ), .Y(n3024) );
  NAND2X1 U3579 ( .A(n3031), .B(n3030), .Y(n2997) );
  NOR2X1 U3580 ( .A(n3029), .B(n3028), .Y(n3031) );
  MXI2X1 U3581 ( .A(n1504), .B(n3027), .S0(n3184), .Y(n3030) );
  NOR2X1 U3582 ( .A(n3212), .B(\R[1][29] ), .Y(n3029) );
  NAND2X1 U3583 ( .A(n3036), .B(n3035), .Y(n2989) );
  NOR2X1 U3584 ( .A(n3034), .B(n3033), .Y(n3036) );
  MXI2X1 U3585 ( .A(n1505), .B(n3032), .S0(n3184), .Y(n3035) );
  NOR2X1 U3586 ( .A(n3213), .B(\R[1][28] ), .Y(n3034) );
  NAND2X1 U3587 ( .A(n3041), .B(n3040), .Y(n2981) );
  NOR2X1 U3588 ( .A(n3039), .B(n3038), .Y(n3041) );
  MXI2X1 U3589 ( .A(n1506), .B(n3037), .S0(n3183), .Y(n3040) );
  NOR2X1 U3590 ( .A(n3206), .B(\R[1][27] ), .Y(n3039) );
  NAND2X1 U3591 ( .A(n3046), .B(n3045), .Y(n2973) );
  NOR2X1 U3592 ( .A(n3044), .B(n3043), .Y(n3046) );
  MXI2X1 U3593 ( .A(n1507), .B(n3042), .S0(n3183), .Y(n3045) );
  NOR2X1 U3594 ( .A(n3213), .B(\R[1][26] ), .Y(n3044) );
  NAND2X1 U3595 ( .A(n3051), .B(n3050), .Y(n2965) );
  NOR2X1 U3596 ( .A(n3049), .B(n3048), .Y(n3051) );
  MXI2X1 U3597 ( .A(n1508), .B(n3047), .S0(n3183), .Y(n3050) );
  NOR2X1 U3598 ( .A(n3210), .B(\R[1][25] ), .Y(n3049) );
  NAND2X1 U3599 ( .A(n3061), .B(n3060), .Y(n2949) );
  NOR2X1 U3600 ( .A(n3059), .B(n3058), .Y(n3061) );
  MXI2X1 U3601 ( .A(n1510), .B(n3057), .S0(n3183), .Y(n3060) );
  NOR2X1 U3602 ( .A(n3210), .B(\R[1][23] ), .Y(n3059) );
  NAND2X1 U3603 ( .A(n3091), .B(n3090), .Y(n2901) );
  NOR2X1 U3604 ( .A(n3089), .B(n3088), .Y(n3091) );
  MXI2X1 U3605 ( .A(n1516), .B(n3087), .S0(n3183), .Y(n3090) );
  NOR2X1 U3606 ( .A(n3211), .B(\R[1][17] ), .Y(n3089) );
  NAND2X1 U3607 ( .A(n3106), .B(n3105), .Y(n2877) );
  NOR2X1 U3608 ( .A(n3104), .B(n3103), .Y(n3106) );
  MXI2X1 U3609 ( .A(n1519), .B(n3102), .S0(n3183), .Y(n3105) );
  NOR2X1 U3610 ( .A(n3211), .B(\R[1][14] ), .Y(n3104) );
  NAND2X1 U3611 ( .A(n3111), .B(n3110), .Y(n2869) );
  NOR2X1 U3612 ( .A(n3109), .B(n3108), .Y(n3111) );
  MXI2X1 U3613 ( .A(n1520), .B(n3107), .S0(n3183), .Y(n3110) );
  NOR2X1 U3614 ( .A(n3211), .B(\R[1][13] ), .Y(n3109) );
  NAND2X1 U3615 ( .A(n3116), .B(n3115), .Y(n2861) );
  NOR2X1 U3616 ( .A(n3114), .B(n3113), .Y(n3116) );
  MXI2X1 U3617 ( .A(n1521), .B(n3112), .S0(n3183), .Y(n3115) );
  NOR2X1 U3618 ( .A(n3212), .B(\R[1][12] ), .Y(n3114) );
  NAND2X1 U3619 ( .A(n3121), .B(n3120), .Y(n2853) );
  NOR2X1 U3620 ( .A(n3119), .B(n3118), .Y(n3121) );
  MXI2X1 U3621 ( .A(n1522), .B(n3117), .S0(n3183), .Y(n3120) );
  NOR2X1 U3622 ( .A(n3212), .B(\R[1][11] ), .Y(n3119) );
  NAND2X1 U3623 ( .A(n3126), .B(n3125), .Y(n2845) );
  NOR2X1 U3624 ( .A(n3124), .B(n3123), .Y(n3126) );
  MXI2X1 U3625 ( .A(n1523), .B(n3122), .S0(n3183), .Y(n3125) );
  NOR2X1 U3626 ( .A(n3212), .B(\R[1][10] ), .Y(n3124) );
  CLKINVX1 U3627 ( .A(instruction[31]), .Y(n3994) );
  MXI4X1 U3628 ( .A(n3381), .B(n3382), .C(n3383), .D(n3384), .S0(n3762), .S1(
        n3754), .Y(n3380) );
  MXI4X1 U3629 ( .A(n3376), .B(n3377), .C(n3378), .D(n3379), .S0(n3762), .S1(
        n3754), .Y(n3375) );
  MXI4X1 U3630 ( .A(\R[12][14] ), .B(\R[13][14] ), .C(\R[14][14] ), .D(
        \R[15][14] ), .S0(n3719), .S1(n3744), .Y(n3384) );
  CLKMX2X2 U3631 ( .A(n3390), .B(n3385), .S0(n3768), .Y(N238) );
  MXI4X1 U3632 ( .A(n3391), .B(n3392), .C(n3393), .D(n3394), .S0(n3762), .S1(
        n3754), .Y(n3390) );
  MXI4X1 U3633 ( .A(n3386), .B(n3387), .C(n3388), .D(n3389), .S0(n3762), .S1(
        n3754), .Y(n3385) );
  MXI4X1 U3634 ( .A(\R[12][15] ), .B(\R[13][15] ), .C(\R[14][15] ), .D(
        \R[15][15] ), .S0(n3719), .S1(n3744), .Y(n3394) );
  CLKMX2X2 U3635 ( .A(n3410), .B(n3405), .S0(n3768), .Y(N236) );
  MXI4X1 U3636 ( .A(n3411), .B(n3412), .C(n3413), .D(n3414), .S0(n3762), .S1(
        n3754), .Y(n3410) );
  MXI4X1 U3637 ( .A(n3406), .B(n3407), .C(n3408), .D(n3409), .S0(n3762), .S1(
        n3754), .Y(n3405) );
  MXI4X1 U3638 ( .A(\R[12][17] ), .B(\R[13][17] ), .C(\R[14][17] ), .D(
        \R[15][17] ), .S0(n3715), .S1(n3744), .Y(n3414) );
  CLKMX2X2 U3639 ( .A(n3400), .B(n3395), .S0(n3768), .Y(N237) );
  MXI4X1 U3640 ( .A(n3401), .B(n3402), .C(n3403), .D(n3404), .S0(n3762), .S1(
        n3754), .Y(n3400) );
  MXI4X1 U3641 ( .A(n3396), .B(n3397), .C(n3398), .D(n3399), .S0(n3762), .S1(
        n3754), .Y(n3395) );
  MXI4X1 U3642 ( .A(\R[12][16] ), .B(\R[13][16] ), .C(\R[14][16] ), .D(
        \R[15][16] ), .S0(n3715), .S1(n3744), .Y(n3404) );
  CLKMX2X2 U3643 ( .A(n3370), .B(n3365), .S0(n3768), .Y(N240) );
  MXI4X1 U3644 ( .A(n3371), .B(n3372), .C(n3373), .D(n3374), .S0(n3761), .S1(
        n3753), .Y(n3370) );
  MXI4X1 U3645 ( .A(n3366), .B(n3367), .C(n3368), .D(n3369), .S0(n3761), .S1(
        n3753), .Y(n3365) );
  MXI4X1 U3646 ( .A(\R[12][13] ), .B(\R[13][13] ), .C(\R[14][13] ), .D(
        \R[15][13] ), .S0(n3718), .S1(n3744), .Y(n3374) );
  OAI22XL U3647 ( .A0(n3899), .A1(n168), .B0(n586), .B1(n3852), .Y(n1620) );
  OAI22XL U3648 ( .A0(n3896), .A1(n168), .B0(n587), .B1(n3852), .Y(n1621) );
  OAI22XL U3649 ( .A0(n3893), .A1(n168), .B0(n588), .B1(n3852), .Y(n1622) );
  OAI22XL U3650 ( .A0(n3890), .A1(n168), .B0(n589), .B1(n3852), .Y(n1623) );
  OAI22XL U3651 ( .A0(n3887), .A1(n168), .B0(n590), .B1(n3852), .Y(n1624) );
  OAI22XL U3652 ( .A0(n3884), .A1(n3851), .B0(n591), .B1(n3852), .Y(n1625) );
  OAI22XL U3653 ( .A0(n3899), .A1(n171), .B0(n618), .B1(n3850), .Y(n1652) );
  OAI22XL U3654 ( .A0(n3896), .A1(n171), .B0(n619), .B1(n3850), .Y(n1653) );
  OAI22XL U3655 ( .A0(n3893), .A1(n171), .B0(n620), .B1(n3850), .Y(n1654) );
  OAI22XL U3656 ( .A0(n3890), .A1(n171), .B0(n621), .B1(n3850), .Y(n1655) );
  OAI22XL U3657 ( .A0(n3887), .A1(n171), .B0(n622), .B1(n3850), .Y(n1656) );
  OAI22XL U3658 ( .A0(n3884), .A1(n3849), .B0(n623), .B1(n3850), .Y(n1657) );
  OAI22XL U3659 ( .A0(n3899), .A1(n175), .B0(n650), .B1(n3845), .Y(n1684) );
  OAI22XL U3660 ( .A0(n3896), .A1(n175), .B0(n651), .B1(n3845), .Y(n1685) );
  OAI22XL U3661 ( .A0(n3893), .A1(n175), .B0(n652), .B1(n3845), .Y(n1686) );
  OAI22XL U3662 ( .A0(n3890), .A1(n175), .B0(n653), .B1(n3845), .Y(n1687) );
  OAI22XL U3663 ( .A0(n3887), .A1(n175), .B0(n654), .B1(n3845), .Y(n1688) );
  OAI22XL U3664 ( .A0(n3884), .A1(n3844), .B0(n655), .B1(n3845), .Y(n1689) );
  OAI22XL U3665 ( .A0(n3899), .A1(n3842), .B0(n682), .B1(n3843), .Y(n1716) );
  OAI22XL U3666 ( .A0(n3896), .A1(n3841), .B0(n683), .B1(n3843), .Y(n1717) );
  OAI22XL U3667 ( .A0(n3893), .A1(n3842), .B0(n684), .B1(n3843), .Y(n1718) );
  OAI22XL U3668 ( .A0(n3890), .A1(n3841), .B0(n685), .B1(n3843), .Y(n1719) );
  OAI22XL U3669 ( .A0(n3887), .A1(n177), .B0(n686), .B1(n3843), .Y(n1720) );
  OAI22XL U3670 ( .A0(n3884), .A1(n3841), .B0(n687), .B1(n3843), .Y(n1721) );
  OAI22XL U3671 ( .A0(n3900), .A1(n181), .B0(n714), .B1(n3840), .Y(n1748) );
  OAI22XL U3672 ( .A0(n3897), .A1(n181), .B0(n715), .B1(n3840), .Y(n1749) );
  OAI22XL U3673 ( .A0(n3894), .A1(n181), .B0(n716), .B1(n3840), .Y(n1750) );
  OAI22XL U3674 ( .A0(n3891), .A1(n181), .B0(n717), .B1(n3840), .Y(n1751) );
  OAI22XL U3675 ( .A0(n3888), .A1(n181), .B0(n718), .B1(n3840), .Y(n1752) );
  OAI22XL U3676 ( .A0(n3885), .A1(n3839), .B0(n719), .B1(n3840), .Y(n1753) );
  OAI22XL U3677 ( .A0(n3900), .A1(n184), .B0(n746), .B1(n3838), .Y(n1780) );
  OAI22XL U3678 ( .A0(n3897), .A1(n184), .B0(n747), .B1(n3838), .Y(n1781) );
  OAI22XL U3679 ( .A0(n3894), .A1(n184), .B0(n748), .B1(n3838), .Y(n1782) );
  OAI22XL U3680 ( .A0(n3891), .A1(n184), .B0(n749), .B1(n3838), .Y(n1783) );
  OAI22XL U3681 ( .A0(n3888), .A1(n184), .B0(n750), .B1(n3838), .Y(n1784) );
  OAI22XL U3682 ( .A0(n3885), .A1(n3837), .B0(n751), .B1(n3838), .Y(n1785) );
  OAI22XL U3683 ( .A0(n3900), .A1(n186), .B0(n778), .B1(n3836), .Y(n1812) );
  OAI22XL U3684 ( .A0(n3897), .A1(n186), .B0(n779), .B1(n3836), .Y(n1813) );
  OAI22XL U3685 ( .A0(n3894), .A1(n186), .B0(n780), .B1(n3836), .Y(n1814) );
  OAI22XL U3686 ( .A0(n3891), .A1(n186), .B0(n781), .B1(n3836), .Y(n1815) );
  OAI22XL U3687 ( .A0(n3888), .A1(n186), .B0(n782), .B1(n3836), .Y(n1816) );
  OAI22XL U3688 ( .A0(n3885), .A1(n3835), .B0(n783), .B1(n3836), .Y(n1817) );
  OAI22XL U3689 ( .A0(n3900), .A1(n3833), .B0(n810), .B1(n3834), .Y(n1844) );
  OAI22XL U3690 ( .A0(n3897), .A1(n3832), .B0(n811), .B1(n3834), .Y(n1845) );
  OAI22XL U3691 ( .A0(n3894), .A1(n3833), .B0(n812), .B1(n3834), .Y(n1846) );
  OAI22XL U3692 ( .A0(n3891), .A1(n3832), .B0(n813), .B1(n3834), .Y(n1847) );
  OAI22XL U3693 ( .A0(n3888), .A1(n188), .B0(n814), .B1(n3834), .Y(n1848) );
  OAI22XL U3694 ( .A0(n3885), .A1(n3832), .B0(n815), .B1(n3834), .Y(n1849) );
  OAI22XL U3695 ( .A0(n3900), .A1(n191), .B0(n842), .B1(n3831), .Y(n1876) );
  OAI22XL U3696 ( .A0(n3897), .A1(n191), .B0(n843), .B1(n3831), .Y(n1877) );
  OAI22XL U3697 ( .A0(n3894), .A1(n191), .B0(n844), .B1(n3831), .Y(n1878) );
  OAI22XL U3698 ( .A0(n3891), .A1(n191), .B0(n845), .B1(n3831), .Y(n1879) );
  OAI22XL U3699 ( .A0(n3888), .A1(n191), .B0(n846), .B1(n3831), .Y(n1880) );
  OAI22XL U3700 ( .A0(n3885), .A1(n3830), .B0(n847), .B1(n3831), .Y(n1881) );
  OAI22XL U3701 ( .A0(n3900), .A1(n194), .B0(n874), .B1(n3829), .Y(n1908) );
  OAI22XL U3702 ( .A0(n3897), .A1(n194), .B0(n875), .B1(n3829), .Y(n1909) );
  OAI22XL U3703 ( .A0(n3894), .A1(n194), .B0(n876), .B1(n3829), .Y(n1910) );
  OAI22XL U3704 ( .A0(n3891), .A1(n194), .B0(n877), .B1(n3829), .Y(n1911) );
  OAI22XL U3705 ( .A0(n3888), .A1(n194), .B0(n878), .B1(n3829), .Y(n1912) );
  OAI22XL U3706 ( .A0(n3885), .A1(n3828), .B0(n879), .B1(n3829), .Y(n1913) );
  OAI22XL U3707 ( .A0(n3900), .A1(n196), .B0(n906), .B1(n3827), .Y(n1940) );
  OAI22XL U3708 ( .A0(n3897), .A1(n196), .B0(n907), .B1(n3827), .Y(n1941) );
  OAI22XL U3709 ( .A0(n3894), .A1(n196), .B0(n908), .B1(n3827), .Y(n1942) );
  OAI22XL U3710 ( .A0(n3891), .A1(n196), .B0(n909), .B1(n3827), .Y(n1943) );
  OAI22XL U3711 ( .A0(n3888), .A1(n196), .B0(n910), .B1(n3827), .Y(n1944) );
  OAI22XL U3712 ( .A0(n3885), .A1(n3826), .B0(n911), .B1(n3827), .Y(n1945) );
  OAI22XL U3713 ( .A0(n3900), .A1(n3824), .B0(n938), .B1(n3825), .Y(n1972) );
  OAI22XL U3714 ( .A0(n3897), .A1(n3823), .B0(n939), .B1(n3825), .Y(n1973) );
  OAI22XL U3715 ( .A0(n3894), .A1(n3824), .B0(n940), .B1(n3825), .Y(n1974) );
  OAI22XL U3716 ( .A0(n3891), .A1(n3823), .B0(n941), .B1(n3825), .Y(n1975) );
  OAI22XL U3717 ( .A0(n3888), .A1(n198), .B0(n942), .B1(n3825), .Y(n1976) );
  OAI22XL U3718 ( .A0(n3885), .A1(n3823), .B0(n943), .B1(n3825), .Y(n1977) );
  OAI22XL U3719 ( .A0(n3900), .A1(n204), .B0(n970), .B1(n3820), .Y(n2004) );
  OAI22XL U3720 ( .A0(n3897), .A1(n204), .B0(n971), .B1(n3820), .Y(n2005) );
  OAI22XL U3721 ( .A0(n3894), .A1(n204), .B0(n972), .B1(n3820), .Y(n2006) );
  OAI22XL U3722 ( .A0(n3891), .A1(n204), .B0(n973), .B1(n3820), .Y(n2007) );
  OAI22XL U3723 ( .A0(n3888), .A1(n204), .B0(n974), .B1(n3820), .Y(n2008) );
  OAI22XL U3724 ( .A0(n3885), .A1(n3819), .B0(n975), .B1(n3820), .Y(n2009) );
  OAI22XL U3725 ( .A0(n3900), .A1(n207), .B0(n1002), .B1(n3818), .Y(n2036) );
  OAI22XL U3726 ( .A0(n3897), .A1(n207), .B0(n1003), .B1(n3818), .Y(n2037) );
  OAI22XL U3727 ( .A0(n3894), .A1(n207), .B0(n1004), .B1(n3818), .Y(n2038) );
  OAI22XL U3728 ( .A0(n3891), .A1(n207), .B0(n1005), .B1(n3818), .Y(n2039) );
  OAI22XL U3729 ( .A0(n3888), .A1(n207), .B0(n1006), .B1(n3818), .Y(n2040) );
  OAI22XL U3730 ( .A0(n3885), .A1(n3817), .B0(n1007), .B1(n3818), .Y(n2041) );
  OAI22XL U3731 ( .A0(n3900), .A1(n209), .B0(n1034), .B1(n3816), .Y(n2068) );
  OAI22XL U3732 ( .A0(n3897), .A1(n209), .B0(n1035), .B1(n3816), .Y(n2069) );
  OAI22XL U3733 ( .A0(n3894), .A1(n209), .B0(n1036), .B1(n3816), .Y(n2070) );
  OAI22XL U3734 ( .A0(n3891), .A1(n209), .B0(n1037), .B1(n3816), .Y(n2071) );
  OAI22XL U3735 ( .A0(n3888), .A1(n209), .B0(n1038), .B1(n3816), .Y(n2072) );
  OAI22XL U3736 ( .A0(n3885), .A1(n3815), .B0(n1039), .B1(n3816), .Y(n2073) );
  OAI22XL U3737 ( .A0(n3901), .A1(n3813), .B0(n1066), .B1(n3814), .Y(n2100) );
  OAI22XL U3738 ( .A0(n3898), .A1(n3812), .B0(n1067), .B1(n3814), .Y(n2101) );
  OAI22XL U3739 ( .A0(n3895), .A1(n3813), .B0(n1068), .B1(n3814), .Y(n2102) );
  OAI22XL U3740 ( .A0(n3892), .A1(n3812), .B0(n1069), .B1(n3814), .Y(n2103) );
  OAI22XL U3741 ( .A0(n3889), .A1(n211), .B0(n1070), .B1(n3814), .Y(n2104) );
  OAI22XL U3742 ( .A0(n3901), .A1(n214), .B0(n1098), .B1(n3811), .Y(n2132) );
  OAI22XL U3743 ( .A0(n3898), .A1(n214), .B0(n1099), .B1(n3811), .Y(n2133) );
  OAI22XL U3744 ( .A0(n3895), .A1(n214), .B0(n1100), .B1(n3811), .Y(n2134) );
  OAI22XL U3745 ( .A0(n3892), .A1(n214), .B0(n1101), .B1(n3811), .Y(n2135) );
  OAI22XL U3746 ( .A0(n3889), .A1(n214), .B0(n1102), .B1(n3811), .Y(n2136) );
  OAI22XL U3747 ( .A0(n3901), .A1(n217), .B0(n1130), .B1(n3808), .Y(n2164) );
  OAI22XL U3748 ( .A0(n3898), .A1(n217), .B0(n1131), .B1(n3808), .Y(n2165) );
  OAI22XL U3749 ( .A0(n3895), .A1(n217), .B0(n1132), .B1(n3808), .Y(n2166) );
  OAI22XL U3750 ( .A0(n3892), .A1(n217), .B0(n1133), .B1(n3808), .Y(n2167) );
  OAI22XL U3751 ( .A0(n3889), .A1(n217), .B0(n1134), .B1(n3808), .Y(n2168) );
  OAI22XL U3752 ( .A0(n3901), .A1(n219), .B0(n1162), .B1(n3805), .Y(n2196) );
  OAI22XL U3753 ( .A0(n3898), .A1(n219), .B0(n1163), .B1(n3805), .Y(n2197) );
  OAI22XL U3754 ( .A0(n3895), .A1(n219), .B0(n1164), .B1(n3805), .Y(n2198) );
  OAI22XL U3755 ( .A0(n3892), .A1(n219), .B0(n1165), .B1(n3805), .Y(n2199) );
  OAI22XL U3756 ( .A0(n3889), .A1(n219), .B0(n1166), .B1(n3805), .Y(n2200) );
  OAI22XL U3757 ( .A0(n3901), .A1(n222), .B0(n1194), .B1(n3803), .Y(n2228) );
  OAI22XL U3758 ( .A0(n3898), .A1(n222), .B0(n1195), .B1(n3803), .Y(n2229) );
  OAI22XL U3759 ( .A0(n3895), .A1(n222), .B0(n1196), .B1(n3803), .Y(n2230) );
  OAI22XL U3760 ( .A0(n3892), .A1(n222), .B0(n1197), .B1(n3803), .Y(n2231) );
  OAI22XL U3761 ( .A0(n3889), .A1(n222), .B0(n1198), .B1(n3803), .Y(n2232) );
  OAI22XL U3762 ( .A0(n3901), .A1(n225), .B0(n1226), .B1(n3800), .Y(n2260) );
  OAI22XL U3763 ( .A0(n3898), .A1(n225), .B0(n1227), .B1(n3800), .Y(n2261) );
  OAI22XL U3764 ( .A0(n3895), .A1(n225), .B0(n1228), .B1(n3800), .Y(n2262) );
  OAI22XL U3765 ( .A0(n3892), .A1(n225), .B0(n1229), .B1(n3800), .Y(n2263) );
  OAI22XL U3766 ( .A0(n3889), .A1(n225), .B0(n1230), .B1(n3800), .Y(n2264) );
  OAI22XL U3767 ( .A0(n1258), .A1(n3798), .B0(n3901), .B1(n3797), .Y(n2292) );
  OAI22XL U3768 ( .A0(n1259), .A1(n3798), .B0(n3898), .B1(n3797), .Y(n2293) );
  OAI22XL U3769 ( .A0(n1260), .A1(n3798), .B0(n3895), .B1(n3797), .Y(n2294) );
  OAI22XL U3770 ( .A0(n1261), .A1(n3798), .B0(n3892), .B1(n3797), .Y(n2295) );
  OAI22XL U3771 ( .A0(n1262), .A1(n3798), .B0(n3889), .B1(n3797), .Y(n2296) );
  OAI22XL U3772 ( .A0(n1263), .A1(n3798), .B0(n3886), .B1(n3797), .Y(n2297) );
  OAI22XL U3773 ( .A0(n3899), .A1(n114), .B0(n1290), .B1(n3963), .Y(n2324) );
  OAI22XL U3774 ( .A0(n3896), .A1(n114), .B0(n1291), .B1(n3963), .Y(n2325) );
  OAI22XL U3775 ( .A0(n3893), .A1(n114), .B0(n1292), .B1(n3963), .Y(n2326) );
  OAI22XL U3776 ( .A0(n3890), .A1(n114), .B0(n1293), .B1(n3963), .Y(n2327) );
  OAI22XL U3777 ( .A0(n3887), .A1(n114), .B0(n1294), .B1(n3963), .Y(n2328) );
  OAI22XL U3778 ( .A0(n3884), .A1(n3962), .B0(n1295), .B1(n3963), .Y(n2329) );
  OAI22XL U3779 ( .A0(n3899), .A1(n149), .B0(n1322), .B1(n3868), .Y(n2356) );
  OAI22XL U3780 ( .A0(n3896), .A1(n149), .B0(n1323), .B1(n3868), .Y(n2357) );
  OAI22XL U3781 ( .A0(n3893), .A1(n149), .B0(n1324), .B1(n3868), .Y(n2358) );
  OAI22XL U3782 ( .A0(n3890), .A1(n149), .B0(n1325), .B1(n3868), .Y(n2359) );
  OAI22XL U3783 ( .A0(n3887), .A1(n149), .B0(n1326), .B1(n3868), .Y(n2360) );
  OAI22XL U3784 ( .A0(n3884), .A1(n3867), .B0(n1327), .B1(n3868), .Y(n2361) );
  OAI22XL U3785 ( .A0(n3899), .A1(n152), .B0(n1354), .B1(n3866), .Y(n2388) );
  OAI22XL U3786 ( .A0(n3896), .A1(n152), .B0(n1355), .B1(n3866), .Y(n2389) );
  OAI22XL U3787 ( .A0(n3893), .A1(n152), .B0(n1356), .B1(n3866), .Y(n2390) );
  OAI22XL U3788 ( .A0(n3890), .A1(n152), .B0(n1357), .B1(n3866), .Y(n2391) );
  OAI22XL U3789 ( .A0(n3887), .A1(n152), .B0(n1358), .B1(n3866), .Y(n2392) );
  OAI22XL U3790 ( .A0(n3884), .A1(n3864), .B0(n1359), .B1(n3866), .Y(n2393) );
  OAI22XL U3791 ( .A0(n3899), .A1(n156), .B0(n1386), .B1(n3863), .Y(n2420) );
  OAI22XL U3792 ( .A0(n3896), .A1(n156), .B0(n1387), .B1(n3863), .Y(n2421) );
  OAI22XL U3793 ( .A0(n3893), .A1(n156), .B0(n1388), .B1(n3863), .Y(n2422) );
  OAI22XL U3794 ( .A0(n3890), .A1(n156), .B0(n1389), .B1(n3863), .Y(n2423) );
  OAI22XL U3795 ( .A0(n3887), .A1(n156), .B0(n1390), .B1(n3863), .Y(n2424) );
  OAI22XL U3796 ( .A0(n3884), .A1(n3861), .B0(n1391), .B1(n3863), .Y(n2425) );
  OAI22XL U3797 ( .A0(n3899), .A1(n159), .B0(n1418), .B1(n3860), .Y(n2452) );
  OAI22XL U3798 ( .A0(n3896), .A1(n159), .B0(n1419), .B1(n3860), .Y(n2453) );
  OAI22XL U3799 ( .A0(n3893), .A1(n159), .B0(n1420), .B1(n3860), .Y(n2454) );
  OAI22XL U3800 ( .A0(n3890), .A1(n159), .B0(n1421), .B1(n3860), .Y(n2455) );
  OAI22XL U3801 ( .A0(n3887), .A1(n159), .B0(n1422), .B1(n3860), .Y(n2456) );
  OAI22XL U3802 ( .A0(n3884), .A1(n3858), .B0(n1423), .B1(n3860), .Y(n2457) );
  OAI22XL U3803 ( .A0(n3899), .A1(n161), .B0(n1450), .B1(n3857), .Y(n2484) );
  OAI22XL U3804 ( .A0(n3896), .A1(n161), .B0(n1451), .B1(n3857), .Y(n2485) );
  OAI22XL U3805 ( .A0(n3893), .A1(n161), .B0(n1452), .B1(n3857), .Y(n2486) );
  OAI22XL U3806 ( .A0(n3890), .A1(n161), .B0(n1453), .B1(n3857), .Y(n2487) );
  OAI22XL U3807 ( .A0(n3887), .A1(n161), .B0(n1454), .B1(n3857), .Y(n2488) );
  OAI22XL U3808 ( .A0(n3884), .A1(n3855), .B0(n1455), .B1(n3857), .Y(n2489) );
  OAI22XL U3809 ( .A0(n3899), .A1(n165), .B0(n1482), .B1(n3854), .Y(n2516) );
  OAI22XL U3810 ( .A0(n3896), .A1(n165), .B0(n1483), .B1(n3854), .Y(n2517) );
  OAI22XL U3811 ( .A0(n3893), .A1(n165), .B0(n1484), .B1(n3854), .Y(n2518) );
  OAI22XL U3812 ( .A0(n3890), .A1(n165), .B0(n1485), .B1(n3854), .Y(n2519) );
  OAI22XL U3813 ( .A0(n3887), .A1(n165), .B0(n1486), .B1(n3854), .Y(n2520) );
  OAI22XL U3814 ( .A0(n3884), .A1(n3853), .B0(n1487), .B1(n3854), .Y(n2521) );
  OAI22XL U3815 ( .A0(n3899), .A1(n3846), .B0(n1514), .B1(n3848), .Y(n2548) );
  OAI22XL U3816 ( .A0(n3896), .A1(n3847), .B0(n1515), .B1(n3848), .Y(n2549) );
  OAI22XL U3817 ( .A0(n3893), .A1(n3846), .B0(n1516), .B1(n3848), .Y(n2550) );
  OAI22XL U3818 ( .A0(n3890), .A1(n173), .B0(n1517), .B1(n3848), .Y(n2551) );
  OAI22XL U3819 ( .A0(n3887), .A1(n173), .B0(n1518), .B1(n3848), .Y(n2552) );
  OAI22XL U3820 ( .A0(n3884), .A1(n3846), .B0(n1519), .B1(n3848), .Y(n2553) );
  OAI22XL U3821 ( .A0(n3900), .A1(n201), .B0(n1546), .B1(n3822), .Y(n2580) );
  OAI22XL U3822 ( .A0(n3897), .A1(n201), .B0(n1547), .B1(n3822), .Y(n2581) );
  OAI22XL U3823 ( .A0(n3894), .A1(n201), .B0(n1548), .B1(n3822), .Y(n2582) );
  OAI22XL U3824 ( .A0(n3891), .A1(n201), .B0(n1549), .B1(n3822), .Y(n2583) );
  OAI22XL U3825 ( .A0(n3888), .A1(n201), .B0(n1550), .B1(n3822), .Y(n2584) );
  OAI22XL U3826 ( .A0(n3885), .A1(n3821), .B0(n1551), .B1(n3822), .Y(n2585) );
  CLKINVX1 U3827 ( .A(instruction[30]), .Y(n3999) );
  AND4X1 U3828 ( .A(n393), .B(n394), .C(n395), .D(n396), .Y(n136) );
  AOI222XL U3829 ( .A0(dataout[19]), .A1(n3771), .B0(N947), .B1(n3775), .C0(
        n3997), .C1(n4013), .Y(n393) );
  AOI222XL U3830 ( .A0(N915), .A1(n253), .B0(N883), .B1(n3778), .C0(N804), 
        .C1(n249), .Y(n394) );
  AOI222XL U3831 ( .A0(N676), .A1(n247), .B0(n2649), .B1(n397), .C0(N234), 
        .C1(n398), .Y(n396) );
  AND4X1 U3832 ( .A(n399), .B(n400), .C(n401), .D(n402), .Y(n137) );
  AOI222XL U3833 ( .A0(dataout[18]), .A1(n3772), .B0(N946), .B1(n3776), .C0(
        n3997), .C1(n2710), .Y(n399) );
  AOI222XL U3834 ( .A0(N914), .A1(n3777), .B0(N882), .B1(n251), .C0(N803), 
        .C1(n3782), .Y(n400) );
  AOI222XL U3835 ( .A0(N675), .A1(n3781), .B0(N203), .B1(n403), .C0(N235), 
        .C1(n404), .Y(n402) );
  AND4X1 U3836 ( .A(n405), .B(n406), .C(n407), .D(n408), .Y(n138) );
  AOI222XL U3837 ( .A0(dataout[17]), .A1(n252), .B0(N945), .B1(n254), .C0(
        n3997), .C1(n2716), .Y(n405) );
  AOI222XL U3838 ( .A0(N913), .A1(n253), .B0(N881), .B1(n3778), .C0(N802), 
        .C1(n249), .Y(n406) );
  AOI222XL U3839 ( .A0(N674), .A1(n247), .B0(N204), .B1(n409), .C0(N236), .C1(
        n410), .Y(n408) );
  AND4X1 U3840 ( .A(n411), .B(n412), .C(n413), .D(n414), .Y(n139) );
  AOI222XL U3841 ( .A0(dataout[16]), .A1(n3771), .B0(N944), .B1(n3775), .C0(
        n3997), .C1(n2713), .Y(n411) );
  AOI222XL U3842 ( .A0(N673), .A1(n3781), .B0(N205), .B1(n415), .C0(N237), 
        .C1(n416), .Y(n414) );
  AOI222XL U3843 ( .A0(N912), .A1(n3777), .B0(N880), .B1(n251), .C0(N801), 
        .C1(n3782), .Y(n412) );
  AND4X1 U3844 ( .A(n417), .B(n418), .C(n419), .D(n420), .Y(n140) );
  AOI222XL U3845 ( .A0(dataout[15]), .A1(n3772), .B0(N943), .B1(n3776), .C0(
        n3997), .C1(n4014), .Y(n417) );
  AOI222XL U3846 ( .A0(N672), .A1(n247), .B0(n2653), .B1(n421), .C0(N238), 
        .C1(n422), .Y(n420) );
  AOI222XL U3847 ( .A0(N911), .A1(n253), .B0(N879), .B1(n3778), .C0(N800), 
        .C1(n249), .Y(n418) );
  AND4X1 U3848 ( .A(n423), .B(n424), .C(n425), .D(n426), .Y(n141) );
  AOI221XL U3849 ( .A0(n427), .A1(n2750), .B0(N207), .B1(n428), .C0(n429), .Y(
        n426) );
  AOI222XL U3850 ( .A0(dataout[14]), .A1(n252), .B0(N910), .B1(n253), .C0(N942), .C1(n3775), .Y(n423) );
  AOI222XL U3851 ( .A0(N799), .A1(n249), .B0(N415), .B1(n250), .C0(N878), .C1(
        n251), .Y(n424) );
  NOR2X1 U3852 ( .A(\R[3][14] ), .B(n3731), .Y(n3640) );
  NOR2X1 U3853 ( .A(\R[3][13] ), .B(n3731), .Y(n3645) );
  NOR2X1 U3854 ( .A(\R[3][17] ), .B(n3730), .Y(n3625) );
  NOR2X1 U3855 ( .A(\R[3][16] ), .B(n3731), .Y(n3630) );
  NOR2X1 U3856 ( .A(\R[3][15] ), .B(n3731), .Y(n3635) );
  NOR2X1 U3857 ( .A(n3748), .B(\R[1][14] ), .Y(n3642) );
  NOR2X1 U3858 ( .A(n3748), .B(\R[1][13] ), .Y(n3647) );
  NOR2X1 U3859 ( .A(n3748), .B(\R[1][16] ), .Y(n3632) );
  NOR2X1 U3860 ( .A(n3748), .B(\R[1][15] ), .Y(n3637) );
  CLKMX2X2 U3861 ( .A(n3360), .B(n3355), .S0(n3768), .Y(N241) );
  MXI4X1 U3862 ( .A(n3361), .B(n3362), .C(n3363), .D(n3364), .S0(n3761), .S1(
        n3753), .Y(n3360) );
  MXI4X1 U3863 ( .A(n3356), .B(n3357), .C(n3358), .D(n3359), .S0(n3761), .S1(
        n3753), .Y(n3355) );
  MXI4X1 U3864 ( .A(\R[12][12] ), .B(\R[13][12] ), .C(\R[14][12] ), .D(
        \R[15][12] ), .S0(n3718), .S1(n3743), .Y(n3364) );
  CLKINVX1 U3865 ( .A(instruction[28]), .Y(n4001) );
  MXI4X1 U3866 ( .A(\R[20][14] ), .B(\R[21][14] ), .C(\R[22][14] ), .D(
        \R[23][14] ), .S0(n3719), .S1(n3744), .Y(n3378) );
  MXI4X1 U3867 ( .A(\R[4][14] ), .B(\R[5][14] ), .C(\R[6][14] ), .D(\R[7][14] ), .S0(n3719), .S1(n3744), .Y(n3383) );
  MXI4X1 U3868 ( .A(\R[20][13] ), .B(\R[21][13] ), .C(\R[22][13] ), .D(
        \R[23][13] ), .S0(n3718), .S1(n3744), .Y(n3368) );
  MXI4X1 U3869 ( .A(\R[4][13] ), .B(\R[5][13] ), .C(\R[6][13] ), .D(\R[7][13] ), .S0(n3719), .S1(n3744), .Y(n3373) );
  MXI4X1 U3870 ( .A(\R[20][15] ), .B(\R[21][15] ), .C(\R[22][15] ), .D(
        \R[23][15] ), .S0(n3719), .S1(n3744), .Y(n3388) );
  MXI4X1 U3871 ( .A(\R[4][15] ), .B(\R[5][15] ), .C(\R[6][15] ), .D(\R[7][15] ), .S0(n3718), .S1(n3744), .Y(n3393) );
  MXI4X1 U3872 ( .A(\R[20][16] ), .B(\R[21][16] ), .C(\R[22][16] ), .D(
        \R[23][16] ), .S0(n3715), .S1(n3744), .Y(n3398) );
  MXI4X1 U3873 ( .A(\R[4][16] ), .B(\R[5][16] ), .C(\R[6][16] ), .D(\R[7][16] ), .S0(n3715), .S1(n3744), .Y(n3403) );
  MXI4X1 U3874 ( .A(\R[16][14] ), .B(\R[17][14] ), .C(\R[18][14] ), .D(
        \R[19][14] ), .S0(n3719), .S1(n3744), .Y(n3376) );
  MXI4X1 U3875 ( .A(\R[16][13] ), .B(\R[17][13] ), .C(\R[18][13] ), .D(
        \R[19][13] ), .S0(n3718), .S1(n3744), .Y(n3366) );
  MXI4X1 U3876 ( .A(\R[16][15] ), .B(\R[17][15] ), .C(\R[18][15] ), .D(
        \R[19][15] ), .S0(n3719), .S1(n3744), .Y(n3386) );
  MXI4X1 U3877 ( .A(\R[16][17] ), .B(\R[17][17] ), .C(\R[18][17] ), .D(
        \R[19][17] ), .S0(n3715), .S1(n3744), .Y(n3406) );
  MXI4X1 U3878 ( .A(\R[16][16] ), .B(\R[17][16] ), .C(\R[18][16] ), .D(
        \R[19][16] ), .S0(n3715), .S1(n3744), .Y(n3396) );
  MXI4X1 U3879 ( .A(\R[24][14] ), .B(\R[25][14] ), .C(\R[26][14] ), .D(
        \R[27][14] ), .S0(n3719), .S1(n3744), .Y(n3377) );
  MXI4X1 U3880 ( .A(\R[8][14] ), .B(\R[9][14] ), .C(\R[10][14] ), .D(
        \R[11][14] ), .S0(n3719), .S1(n3744), .Y(n3382) );
  MXI4X1 U3881 ( .A(\R[24][13] ), .B(\R[25][13] ), .C(\R[26][13] ), .D(
        \R[27][13] ), .S0(n3718), .S1(n3743), .Y(n3367) );
  MXI4X1 U3882 ( .A(\R[8][13] ), .B(\R[9][13] ), .C(\R[10][13] ), .D(
        \R[11][13] ), .S0(n3718), .S1(n3744), .Y(n3372) );
  MXI4X1 U3883 ( .A(\R[24][15] ), .B(\R[25][15] ), .C(\R[26][15] ), .D(
        \R[27][15] ), .S0(n3719), .S1(n3744), .Y(n3387) );
  MXI4X1 U3884 ( .A(\R[8][15] ), .B(\R[9][15] ), .C(\R[10][15] ), .D(
        \R[11][15] ), .S0(n3719), .S1(n3744), .Y(n3392) );
  MXI4X1 U3885 ( .A(\R[24][17] ), .B(\R[25][17] ), .C(\R[26][17] ), .D(
        \R[27][17] ), .S0(n3715), .S1(n3744), .Y(n3407) );
  MXI4X1 U3886 ( .A(\R[24][16] ), .B(\R[25][16] ), .C(\R[26][16] ), .D(
        \R[27][16] ), .S0(n3715), .S1(n3744), .Y(n3397) );
  MXI4X1 U3887 ( .A(\R[8][16] ), .B(\R[9][16] ), .C(\R[10][16] ), .D(
        \R[11][16] ), .S0(n3715), .S1(n3744), .Y(n3402) );
  MXI4X1 U3888 ( .A(\R[28][14] ), .B(\R[29][14] ), .C(\R[30][14] ), .D(
        \R[31][14] ), .S0(n3719), .S1(n3744), .Y(n3379) );
  MXI4X1 U3889 ( .A(\R[28][13] ), .B(\R[29][13] ), .C(\R[30][13] ), .D(
        \R[31][13] ), .S0(n3718), .S1(n3743), .Y(n3369) );
  MXI4X1 U3890 ( .A(\R[28][15] ), .B(\R[29][15] ), .C(\R[30][15] ), .D(
        \R[31][15] ), .S0(n3719), .S1(n3744), .Y(n3389) );
  MXI4X1 U3891 ( .A(\R[28][16] ), .B(\R[29][16] ), .C(\R[30][16] ), .D(
        \R[31][16] ), .S0(n3715), .S1(n3744), .Y(n3399) );
  CLKBUFX3 U3892 ( .A(N48), .Y(n3222) );
  CLKBUFX3 U3893 ( .A(N48), .Y(n3221) );
  CLKBUFX3 U3894 ( .A(N50), .Y(n3234) );
  OAI221XL U3895 ( .A0(n4010), .A1(n3783), .B0(n1568), .B1(n4045), .C0(n493), 
        .Y(n2602) );
  OAI221XL U3896 ( .A0(n2704), .A1(n478), .B0(n1569), .B1(n4045), .C0(n494), 
        .Y(n2603) );
  OAI221XL U3897 ( .A0(n4011), .A1(n3783), .B0(n1570), .B1(n4045), .C0(n495), 
        .Y(n2604) );
  OAI221XL U3898 ( .A0(n2699), .A1(n478), .B0(n1571), .B1(n4045), .C0(n496), 
        .Y(n2605) );
  OAI221XL U3899 ( .A0(n2725), .A1(n3783), .B0(n1572), .B1(n4045), .C0(n497), 
        .Y(n2606) );
  AOI22X1 U3900 ( .A0(N277), .A1(n3789), .B0(N1016), .B1(n3785), .Y(n497) );
  OAI221XL U3901 ( .A0(n2707), .A1(n478), .B0(n1573), .B1(n4045), .C0(n498), 
        .Y(n2607) );
  AOI22X1 U3902 ( .A0(N276), .A1(n3789), .B0(N1015), .B1(n3785), .Y(n498) );
  AND2X2 U3903 ( .A(N91), .B(n3973), .Y(N157) );
  CLKMX2X2 U3904 ( .A(n3450), .B(n3445), .S0(n3769), .Y(N232) );
  MXI4X1 U3905 ( .A(n3451), .B(n3452), .C(n3453), .D(n3454), .S0(n3763), .S1(
        n3755), .Y(n3450) );
  MXI4X1 U3906 ( .A(n3446), .B(n3447), .C(n3448), .D(n3449), .S0(n3763), .S1(
        n3755), .Y(n3445) );
  MXI4X1 U3907 ( .A(\R[12][21] ), .B(\R[13][21] ), .C(\R[14][21] ), .D(
        \R[15][21] ), .S0(n3716), .S1(n3744), .Y(n3454) );
  CLKMX2X2 U3908 ( .A(n3430), .B(n3425), .S0(n3768), .Y(N234) );
  MXI4X1 U3909 ( .A(n3431), .B(n3432), .C(n3433), .D(n3434), .S0(n3762), .S1(
        n3754), .Y(n3430) );
  MXI4X1 U3910 ( .A(n3426), .B(n3427), .C(n3428), .D(n3429), .S0(n3762), .S1(
        n3754), .Y(n3425) );
  MXI4X1 U3911 ( .A(\R[12][19] ), .B(\R[13][19] ), .C(\R[14][19] ), .D(
        \R[15][19] ), .S0(n3715), .S1(n3744), .Y(n3434) );
  CLKMX2X2 U3912 ( .A(n3460), .B(n3455), .S0(n3769), .Y(N231) );
  MXI4X1 U3913 ( .A(n3461), .B(n3462), .C(n3463), .D(n3464), .S0(n3763), .S1(
        n3755), .Y(n3460) );
  MXI4X1 U3914 ( .A(n3456), .B(n3457), .C(n3458), .D(n3459), .S0(n3763), .S1(
        n3755), .Y(n3455) );
  MXI4X1 U3915 ( .A(\R[12][22] ), .B(\R[13][22] ), .C(\R[14][22] ), .D(
        \R[15][22] ), .S0(n3716), .S1(n3745), .Y(n3464) );
  CLKMX2X2 U3916 ( .A(n3440), .B(n3435), .S0(n3769), .Y(N233) );
  MXI4X1 U3917 ( .A(n3441), .B(n3442), .C(n3443), .D(n3444), .S0(n3763), .S1(
        n3755), .Y(n3440) );
  MXI4X1 U3918 ( .A(n3436), .B(n3437), .C(n3438), .D(n3439), .S0(n3763), .S1(
        n3755), .Y(n3435) );
  MXI4X1 U3919 ( .A(\R[12][20] ), .B(\R[13][20] ), .C(\R[14][20] ), .D(
        \R[15][20] ), .S0(n3715), .S1(n3744), .Y(n3444) );
  CLKMX2X2 U3920 ( .A(n3420), .B(n3415), .S0(n3768), .Y(N235) );
  MXI4X1 U3921 ( .A(n3421), .B(n3422), .C(n3423), .D(n3424), .S0(n3762), .S1(
        n3754), .Y(n3420) );
  MXI4X1 U3922 ( .A(n3416), .B(n3417), .C(n3418), .D(n3419), .S0(n3762), .S1(
        n3754), .Y(n3415) );
  MXI4X1 U3923 ( .A(\R[12][18] ), .B(\R[13][18] ), .C(\R[14][18] ), .D(
        \R[15][18] ), .S0(n3715), .S1(n3744), .Y(n3424) );
  OAI22XL U3924 ( .A0(n3881), .A1(n3851), .B0(n592), .B1(n3852), .Y(n1626) );
  OAI22XL U3925 ( .A0(n3878), .A1(n3851), .B0(n593), .B1(n3852), .Y(n1627) );
  OAI22XL U3926 ( .A0(n3875), .A1(n3851), .B0(n594), .B1(n3852), .Y(n1628) );
  OAI22XL U3927 ( .A0(n3872), .A1(n3851), .B0(n595), .B1(n3852), .Y(n1629) );
  OAI22XL U3928 ( .A0(n3964), .A1(n168), .B0(n596), .B1(n3852), .Y(n1630) );
  OAI22XL U3929 ( .A0(n3944), .A1(n168), .B0(n602), .B1(n3852), .Y(n1636) );
  OAI22XL U3930 ( .A0(n3881), .A1(n3849), .B0(n624), .B1(n3850), .Y(n1658) );
  OAI22XL U3931 ( .A0(n3878), .A1(n3849), .B0(n625), .B1(n3850), .Y(n1659) );
  OAI22XL U3932 ( .A0(n3875), .A1(n3849), .B0(n626), .B1(n3850), .Y(n1660) );
  OAI22XL U3933 ( .A0(n3872), .A1(n3849), .B0(n627), .B1(n3850), .Y(n1661) );
  OAI22XL U3934 ( .A0(n3964), .A1(n3849), .B0(n628), .B1(n3850), .Y(n1662) );
  OAI22XL U3935 ( .A0(n3944), .A1(n3849), .B0(n634), .B1(n3850), .Y(n1668) );
  OAI22XL U3936 ( .A0(n3881), .A1(n3844), .B0(n656), .B1(n3845), .Y(n1690) );
  OAI22XL U3937 ( .A0(n3878), .A1(n3844), .B0(n657), .B1(n3845), .Y(n1691) );
  OAI22XL U3938 ( .A0(n3875), .A1(n3844), .B0(n658), .B1(n3845), .Y(n1692) );
  OAI22XL U3939 ( .A0(n3872), .A1(n3844), .B0(n659), .B1(n3845), .Y(n1693) );
  OAI22XL U3940 ( .A0(n3964), .A1(n175), .B0(n660), .B1(n3845), .Y(n1694) );
  OAI22XL U3941 ( .A0(n3944), .A1(n175), .B0(n666), .B1(n3845), .Y(n1700) );
  OAI22XL U3942 ( .A0(n3881), .A1(n3841), .B0(n688), .B1(n3843), .Y(n1722) );
  OAI22XL U3943 ( .A0(n3878), .A1(n3841), .B0(n689), .B1(n3843), .Y(n1723) );
  OAI22XL U3944 ( .A0(n3875), .A1(n3841), .B0(n690), .B1(n3843), .Y(n1724) );
  OAI22XL U3945 ( .A0(n3872), .A1(n3842), .B0(n691), .B1(n3843), .Y(n1725) );
  OAI22XL U3946 ( .A0(n3964), .A1(n3841), .B0(n692), .B1(n3843), .Y(n1726) );
  OAI22XL U3947 ( .A0(n3944), .A1(n3842), .B0(n698), .B1(n3843), .Y(n1732) );
  OAI22XL U3948 ( .A0(n3882), .A1(n3839), .B0(n720), .B1(n3840), .Y(n1754) );
  OAI22XL U3949 ( .A0(n3879), .A1(n3839), .B0(n721), .B1(n3840), .Y(n1755) );
  OAI22XL U3950 ( .A0(n3876), .A1(n3839), .B0(n722), .B1(n3840), .Y(n1756) );
  OAI22XL U3951 ( .A0(n3873), .A1(n3839), .B0(n723), .B1(n3840), .Y(n1757) );
  OAI22XL U3952 ( .A0(n3965), .A1(n3839), .B0(n724), .B1(n3840), .Y(n1758) );
  OAI22XL U3953 ( .A0(n3945), .A1(n3839), .B0(n730), .B1(n3840), .Y(n1764) );
  OAI22XL U3954 ( .A0(n3882), .A1(n3837), .B0(n752), .B1(n3838), .Y(n1786) );
  OAI22XL U3955 ( .A0(n3879), .A1(n3837), .B0(n753), .B1(n3838), .Y(n1787) );
  OAI22XL U3956 ( .A0(n3876), .A1(n3837), .B0(n754), .B1(n3838), .Y(n1788) );
  OAI22XL U3957 ( .A0(n3873), .A1(n3837), .B0(n755), .B1(n3838), .Y(n1789) );
  OAI22XL U3958 ( .A0(n3965), .A1(n3837), .B0(n756), .B1(n3838), .Y(n1790) );
  OAI22XL U3959 ( .A0(n3945), .A1(n3837), .B0(n762), .B1(n3838), .Y(n1796) );
  OAI22XL U3960 ( .A0(n3882), .A1(n3835), .B0(n784), .B1(n3836), .Y(n1818) );
  OAI22XL U3961 ( .A0(n3879), .A1(n3835), .B0(n785), .B1(n3836), .Y(n1819) );
  OAI22XL U3962 ( .A0(n3876), .A1(n3835), .B0(n786), .B1(n3836), .Y(n1820) );
  OAI22XL U3963 ( .A0(n3873), .A1(n3835), .B0(n787), .B1(n3836), .Y(n1821) );
  OAI22XL U3964 ( .A0(n3965), .A1(n186), .B0(n788), .B1(n3836), .Y(n1822) );
  OAI22XL U3965 ( .A0(n3945), .A1(n186), .B0(n794), .B1(n3836), .Y(n1828) );
  OAI22XL U3966 ( .A0(n3882), .A1(n3832), .B0(n816), .B1(n3834), .Y(n1850) );
  OAI22XL U3967 ( .A0(n3879), .A1(n3832), .B0(n817), .B1(n3834), .Y(n1851) );
  OAI22XL U3968 ( .A0(n3876), .A1(n3832), .B0(n818), .B1(n3834), .Y(n1852) );
  OAI22XL U3969 ( .A0(n3873), .A1(n3833), .B0(n819), .B1(n3834), .Y(n1853) );
  OAI22XL U3970 ( .A0(n3965), .A1(n3832), .B0(n820), .B1(n3834), .Y(n1854) );
  OAI22XL U3971 ( .A0(n3945), .A1(n3833), .B0(n826), .B1(n3834), .Y(n1860) );
  OAI22XL U3972 ( .A0(n3882), .A1(n3830), .B0(n848), .B1(n3831), .Y(n1882) );
  OAI22XL U3973 ( .A0(n3879), .A1(n3830), .B0(n849), .B1(n3831), .Y(n1883) );
  OAI22XL U3974 ( .A0(n3876), .A1(n3830), .B0(n850), .B1(n3831), .Y(n1884) );
  OAI22XL U3975 ( .A0(n3873), .A1(n3830), .B0(n851), .B1(n3831), .Y(n1885) );
  OAI22XL U3976 ( .A0(n3965), .A1(n191), .B0(n852), .B1(n3831), .Y(n1886) );
  OAI22XL U3977 ( .A0(n3945), .A1(n191), .B0(n858), .B1(n3831), .Y(n1892) );
  OAI22XL U3978 ( .A0(n3882), .A1(n3828), .B0(n880), .B1(n3829), .Y(n1914) );
  OAI22XL U3979 ( .A0(n3879), .A1(n3828), .B0(n881), .B1(n3829), .Y(n1915) );
  OAI22XL U3980 ( .A0(n3876), .A1(n3828), .B0(n882), .B1(n3829), .Y(n1916) );
  OAI22XL U3981 ( .A0(n3873), .A1(n3828), .B0(n883), .B1(n3829), .Y(n1917) );
  OAI22XL U3982 ( .A0(n3965), .A1(n3828), .B0(n884), .B1(n3829), .Y(n1918) );
  OAI22XL U3983 ( .A0(n3945), .A1(n3828), .B0(n890), .B1(n3829), .Y(n1924) );
  OAI22XL U3984 ( .A0(n3882), .A1(n3826), .B0(n912), .B1(n3827), .Y(n1946) );
  OAI22XL U3985 ( .A0(n3879), .A1(n3826), .B0(n913), .B1(n3827), .Y(n1947) );
  OAI22XL U3986 ( .A0(n3876), .A1(n3826), .B0(n914), .B1(n3827), .Y(n1948) );
  OAI22XL U3987 ( .A0(n3873), .A1(n3826), .B0(n915), .B1(n3827), .Y(n1949) );
  OAI22XL U3988 ( .A0(n3965), .A1(n196), .B0(n916), .B1(n3827), .Y(n1950) );
  OAI22XL U3989 ( .A0(n3945), .A1(n196), .B0(n922), .B1(n3827), .Y(n1956) );
  OAI22XL U3990 ( .A0(n3882), .A1(n3823), .B0(n944), .B1(n3825), .Y(n1978) );
  OAI22XL U3991 ( .A0(n3879), .A1(n3823), .B0(n945), .B1(n3825), .Y(n1979) );
  OAI22XL U3992 ( .A0(n3876), .A1(n3823), .B0(n946), .B1(n3825), .Y(n1980) );
  OAI22XL U3993 ( .A0(n3873), .A1(n3824), .B0(n947), .B1(n3825), .Y(n1981) );
  OAI22XL U3994 ( .A0(n3965), .A1(n3823), .B0(n948), .B1(n3825), .Y(n1982) );
  OAI22XL U3995 ( .A0(n3945), .A1(n3824), .B0(n954), .B1(n3825), .Y(n1988) );
  OAI22XL U3996 ( .A0(n3882), .A1(n3819), .B0(n976), .B1(n3820), .Y(n2010) );
  OAI22XL U3997 ( .A0(n3879), .A1(n3819), .B0(n977), .B1(n3820), .Y(n2011) );
  OAI22XL U3998 ( .A0(n3876), .A1(n3819), .B0(n978), .B1(n3820), .Y(n2012) );
  OAI22XL U3999 ( .A0(n3873), .A1(n3819), .B0(n979), .B1(n3820), .Y(n2013) );
  OAI22XL U4000 ( .A0(n3965), .A1(n204), .B0(n980), .B1(n3820), .Y(n2014) );
  OAI22XL U4001 ( .A0(n3945), .A1(n204), .B0(n986), .B1(n3820), .Y(n2020) );
  OAI22XL U4002 ( .A0(n3882), .A1(n3817), .B0(n1008), .B1(n3818), .Y(n2042) );
  OAI22XL U4003 ( .A0(n3879), .A1(n3817), .B0(n1009), .B1(n3818), .Y(n2043) );
  OAI22XL U4004 ( .A0(n3876), .A1(n3817), .B0(n1010), .B1(n3818), .Y(n2044) );
  OAI22XL U4005 ( .A0(n3873), .A1(n3817), .B0(n1011), .B1(n3818), .Y(n2045) );
  OAI22XL U4006 ( .A0(n3965), .A1(n3817), .B0(n1012), .B1(n3818), .Y(n2046) );
  OAI22XL U4007 ( .A0(n3945), .A1(n3817), .B0(n1018), .B1(n3818), .Y(n2052) );
  OAI22XL U4008 ( .A0(n3882), .A1(n3815), .B0(n1040), .B1(n3816), .Y(n2074) );
  OAI22XL U4009 ( .A0(n3879), .A1(n3815), .B0(n1041), .B1(n3816), .Y(n2075) );
  OAI22XL U4010 ( .A0(n3876), .A1(n3815), .B0(n1042), .B1(n3816), .Y(n2076) );
  OAI22XL U4011 ( .A0(n3873), .A1(n3815), .B0(n1043), .B1(n3816), .Y(n2077) );
  OAI22XL U4012 ( .A0(n3965), .A1(n209), .B0(n1044), .B1(n3816), .Y(n2078) );
  OAI22XL U4013 ( .A0(n3945), .A1(n209), .B0(n1050), .B1(n3816), .Y(n2084) );
  OAI22XL U4014 ( .A0(n3886), .A1(n3812), .B0(n1071), .B1(n3814), .Y(n2105) );
  OAI22XL U4015 ( .A0(n3883), .A1(n3812), .B0(n1072), .B1(n3814), .Y(n2106) );
  OAI22XL U4016 ( .A0(n3880), .A1(n3812), .B0(n1073), .B1(n3814), .Y(n2107) );
  OAI22XL U4017 ( .A0(n3877), .A1(n3812), .B0(n1074), .B1(n3814), .Y(n2108) );
  OAI22XL U4018 ( .A0(n3874), .A1(n3813), .B0(n1075), .B1(n3814), .Y(n2109) );
  OAI22XL U4019 ( .A0(n3966), .A1(n3812), .B0(n1076), .B1(n3814), .Y(n2110) );
  OAI22XL U4020 ( .A0(n3946), .A1(n3813), .B0(n1082), .B1(n3814), .Y(n2116) );
  OAI22XL U4021 ( .A0(n3886), .A1(n3809), .B0(n1103), .B1(n3811), .Y(n2137) );
  OAI22XL U4022 ( .A0(n3883), .A1(n3809), .B0(n1104), .B1(n3811), .Y(n2138) );
  OAI22XL U4023 ( .A0(n3880), .A1(n3809), .B0(n1105), .B1(n3811), .Y(n2139) );
  OAI22XL U4024 ( .A0(n3877), .A1(n3809), .B0(n1106), .B1(n3811), .Y(n2140) );
  OAI22XL U4025 ( .A0(n3874), .A1(n214), .B0(n1107), .B1(n3811), .Y(n2141) );
  OAI22XL U4026 ( .A0(n3966), .A1(n214), .B0(n1108), .B1(n3811), .Y(n2142) );
  OAI22XL U4027 ( .A0(n3946), .A1(n214), .B0(n1114), .B1(n3810), .Y(n2148) );
  OAI22XL U4028 ( .A0(n3886), .A1(n3806), .B0(n1135), .B1(n3808), .Y(n2169) );
  OAI22XL U4029 ( .A0(n3883), .A1(n3806), .B0(n1136), .B1(n3808), .Y(n2170) );
  OAI22XL U4030 ( .A0(n3880), .A1(n3806), .B0(n1137), .B1(n3808), .Y(n2171) );
  OAI22XL U4031 ( .A0(n3877), .A1(n3806), .B0(n1138), .B1(n3808), .Y(n2172) );
  OAI22XL U4032 ( .A0(n3874), .A1(n217), .B0(n1139), .B1(n3808), .Y(n2173) );
  OAI22XL U4033 ( .A0(n3966), .A1(n217), .B0(n1140), .B1(n3808), .Y(n2174) );
  OAI22XL U4034 ( .A0(n3946), .A1(n217), .B0(n1146), .B1(n3807), .Y(n2180) );
  OAI22XL U4035 ( .A0(n3886), .A1(n3804), .B0(n1167), .B1(n3805), .Y(n2201) );
  OAI22XL U4036 ( .A0(n3883), .A1(n3804), .B0(n1168), .B1(n3805), .Y(n2202) );
  OAI22XL U4037 ( .A0(n3880), .A1(n3804), .B0(n1169), .B1(n3805), .Y(n2203) );
  OAI22XL U4038 ( .A0(n3877), .A1(n3804), .B0(n1170), .B1(n3805), .Y(n2204) );
  OAI22XL U4039 ( .A0(n3874), .A1(n3804), .B0(n1171), .B1(n3805), .Y(n2205) );
  OAI22XL U4040 ( .A0(n3966), .A1(n219), .B0(n1172), .B1(n3805), .Y(n2206) );
  OAI22XL U4041 ( .A0(n3946), .A1(n219), .B0(n1178), .B1(n3805), .Y(n2212) );
  OAI22XL U4042 ( .A0(n3886), .A1(n3801), .B0(n1199), .B1(n3803), .Y(n2233) );
  OAI22XL U4043 ( .A0(n3883), .A1(n3801), .B0(n1200), .B1(n3803), .Y(n2234) );
  OAI22XL U4044 ( .A0(n3880), .A1(n3801), .B0(n1201), .B1(n3803), .Y(n2235) );
  OAI22XL U4045 ( .A0(n3877), .A1(n3801), .B0(n1202), .B1(n3803), .Y(n2236) );
  OAI22XL U4046 ( .A0(n3874), .A1(n222), .B0(n1203), .B1(n3803), .Y(n2237) );
  OAI22XL U4047 ( .A0(n3966), .A1(n222), .B0(n1204), .B1(n3803), .Y(n2238) );
  OAI22XL U4048 ( .A0(n3946), .A1(n222), .B0(n1210), .B1(n3802), .Y(n2244) );
  OAI22XL U4049 ( .A0(n3886), .A1(n3799), .B0(n1231), .B1(n3800), .Y(n2265) );
  OAI22XL U4050 ( .A0(n3883), .A1(n3799), .B0(n1232), .B1(n3800), .Y(n2266) );
  OAI22XL U4051 ( .A0(n3880), .A1(n3799), .B0(n1233), .B1(n3800), .Y(n2267) );
  OAI22XL U4052 ( .A0(n3877), .A1(n3799), .B0(n1234), .B1(n3800), .Y(n2268) );
  OAI22XL U4053 ( .A0(n3874), .A1(n3799), .B0(n1235), .B1(n3800), .Y(n2269) );
  OAI22XL U4054 ( .A0(n3966), .A1(n225), .B0(n1236), .B1(n3800), .Y(n2270) );
  OAI22XL U4055 ( .A0(n3946), .A1(n225), .B0(n1242), .B1(n3800), .Y(n2276) );
  OAI22XL U4056 ( .A0(n1264), .A1(n3798), .B0(n3883), .B1(n3797), .Y(n2298) );
  OAI22XL U4057 ( .A0(n1265), .A1(n3798), .B0(n3880), .B1(n3797), .Y(n2299) );
  OAI22XL U4058 ( .A0(n1266), .A1(n3798), .B0(n3877), .B1(n3797), .Y(n2300) );
  OAI22XL U4059 ( .A0(n1267), .A1(n3798), .B0(n3874), .B1(n3795), .Y(n2301) );
  OAI22XL U4060 ( .A0(n1268), .A1(n3798), .B0(n3966), .B1(n3795), .Y(n2302) );
  OAI22XL U4061 ( .A0(n1274), .A1(n3798), .B0(n3946), .B1(n3795), .Y(n2308) );
  OAI22XL U4062 ( .A0(n3881), .A1(n3962), .B0(n1296), .B1(n3963), .Y(n2330) );
  OAI22XL U4063 ( .A0(n3878), .A1(n3962), .B0(n1297), .B1(n3963), .Y(n2331) );
  OAI22XL U4064 ( .A0(n3875), .A1(n3962), .B0(n1298), .B1(n3963), .Y(n2332) );
  OAI22XL U4065 ( .A0(n3872), .A1(n3962), .B0(n1299), .B1(n3963), .Y(n2333) );
  OAI22XL U4066 ( .A0(n3964), .A1(n114), .B0(n1300), .B1(n3963), .Y(n2334) );
  OAI22XL U4067 ( .A0(n3944), .A1(n114), .B0(n1306), .B1(n3963), .Y(n2340) );
  OAI22XL U4068 ( .A0(n3881), .A1(n3867), .B0(n1328), .B1(n3868), .Y(n2362) );
  OAI22XL U4069 ( .A0(n3878), .A1(n3867), .B0(n1329), .B1(n3868), .Y(n2363) );
  OAI22XL U4070 ( .A0(n3875), .A1(n3867), .B0(n1330), .B1(n3868), .Y(n2364) );
  OAI22XL U4071 ( .A0(n3872), .A1(n3867), .B0(n1331), .B1(n3868), .Y(n2365) );
  OAI22XL U4072 ( .A0(n3964), .A1(n149), .B0(n1332), .B1(n3868), .Y(n2366) );
  OAI22XL U4073 ( .A0(n3944), .A1(n149), .B0(n1338), .B1(n3868), .Y(n2372) );
  OAI22XL U4074 ( .A0(n3881), .A1(n3864), .B0(n1360), .B1(n3866), .Y(n2394) );
  OAI22XL U4075 ( .A0(n3878), .A1(n3864), .B0(n1361), .B1(n3866), .Y(n2395) );
  OAI22XL U4076 ( .A0(n3875), .A1(n3864), .B0(n1362), .B1(n3866), .Y(n2396) );
  OAI22XL U4077 ( .A0(n3872), .A1(n3864), .B0(n1363), .B1(n3866), .Y(n2397) );
  OAI22XL U4078 ( .A0(n3964), .A1(n152), .B0(n1364), .B1(n3866), .Y(n2398) );
  OAI22XL U4079 ( .A0(n3944), .A1(n152), .B0(n1370), .B1(n3865), .Y(n2404) );
  OAI22XL U4080 ( .A0(n3881), .A1(n3861), .B0(n1392), .B1(n3863), .Y(n2426) );
  OAI22XL U4081 ( .A0(n3878), .A1(n3861), .B0(n1393), .B1(n3863), .Y(n2427) );
  OAI22XL U4082 ( .A0(n3875), .A1(n3861), .B0(n1394), .B1(n3863), .Y(n2428) );
  OAI22XL U4083 ( .A0(n3872), .A1(n3861), .B0(n1395), .B1(n3863), .Y(n2429) );
  OAI22XL U4084 ( .A0(n3964), .A1(n156), .B0(n1396), .B1(n3863), .Y(n2430) );
  OAI22XL U4085 ( .A0(n3944), .A1(n156), .B0(n1402), .B1(n3862), .Y(n2436) );
  OAI22XL U4086 ( .A0(n3881), .A1(n3858), .B0(n1424), .B1(n3860), .Y(n2458) );
  OAI22XL U4087 ( .A0(n3878), .A1(n3858), .B0(n1425), .B1(n3860), .Y(n2459) );
  OAI22XL U4088 ( .A0(n3875), .A1(n3858), .B0(n1426), .B1(n3860), .Y(n2460) );
  OAI22XL U4089 ( .A0(n3872), .A1(n159), .B0(n1427), .B1(n3860), .Y(n2461) );
  OAI22XL U4090 ( .A0(n3964), .A1(n159), .B0(n1428), .B1(n3860), .Y(n2462) );
  OAI22XL U4091 ( .A0(n3944), .A1(n159), .B0(n1434), .B1(n3859), .Y(n2468) );
  OAI22XL U4092 ( .A0(n3881), .A1(n3855), .B0(n1456), .B1(n3857), .Y(n2490) );
  OAI22XL U4093 ( .A0(n3878), .A1(n3855), .B0(n1457), .B1(n3857), .Y(n2491) );
  OAI22XL U4094 ( .A0(n3875), .A1(n3855), .B0(n1458), .B1(n3857), .Y(n2492) );
  OAI22XL U4095 ( .A0(n3872), .A1(n161), .B0(n1459), .B1(n3857), .Y(n2493) );
  OAI22XL U4096 ( .A0(n3964), .A1(n161), .B0(n1460), .B1(n3857), .Y(n2494) );
  OAI22XL U4097 ( .A0(n3944), .A1(n161), .B0(n1466), .B1(n3856), .Y(n2500) );
  OAI22XL U4098 ( .A0(n3881), .A1(n3853), .B0(n1488), .B1(n3854), .Y(n2522) );
  OAI22XL U4099 ( .A0(n3878), .A1(n3853), .B0(n1489), .B1(n3854), .Y(n2523) );
  OAI22XL U4100 ( .A0(n3875), .A1(n3853), .B0(n1490), .B1(n3854), .Y(n2524) );
  OAI22XL U4101 ( .A0(n3872), .A1(n3853), .B0(n1491), .B1(n3854), .Y(n2525) );
  OAI22XL U4102 ( .A0(n3964), .A1(n165), .B0(n1492), .B1(n3854), .Y(n2526) );
  OAI22XL U4103 ( .A0(n3944), .A1(n165), .B0(n1498), .B1(n3854), .Y(n2532) );
  OAI22XL U4104 ( .A0(n3881), .A1(n3846), .B0(n1520), .B1(n3848), .Y(n2554) );
  OAI22XL U4105 ( .A0(n3878), .A1(n3846), .B0(n1521), .B1(n3848), .Y(n2555) );
  OAI22XL U4106 ( .A0(n3875), .A1(n3846), .B0(n1522), .B1(n3848), .Y(n2556) );
  OAI22XL U4107 ( .A0(n3872), .A1(n3847), .B0(n1523), .B1(n3848), .Y(n2557) );
  OAI22XL U4108 ( .A0(n3964), .A1(n3847), .B0(n1524), .B1(n3848), .Y(n2558) );
  OAI22XL U4109 ( .A0(n3944), .A1(n3847), .B0(n1530), .B1(n3848), .Y(n2564) );
  OAI22XL U4110 ( .A0(n3882), .A1(n3821), .B0(n1552), .B1(n3822), .Y(n2586) );
  OAI22XL U4111 ( .A0(n3879), .A1(n3821), .B0(n1553), .B1(n3822), .Y(n2587) );
  OAI22XL U4112 ( .A0(n3876), .A1(n3821), .B0(n1554), .B1(n3822), .Y(n2588) );
  OAI22XL U4113 ( .A0(n3873), .A1(n3821), .B0(n1555), .B1(n3822), .Y(n2589) );
  OAI22XL U4114 ( .A0(n3965), .A1(n201), .B0(n1556), .B1(n3822), .Y(n2590) );
  OAI22XL U4115 ( .A0(n3945), .A1(n201), .B0(n1562), .B1(n3822), .Y(n2596) );
  AND4X1 U4116 ( .A(n431), .B(n432), .C(n433), .D(n434), .Y(n142) );
  AOI221XL U4117 ( .A0(n435), .A1(n2741), .B0(N208), .B1(n436), .C0(n437), .Y(
        n434) );
  AOI222XL U4118 ( .A0(dataout[13]), .A1(n3771), .B0(N909), .B1(n253), .C0(
        N941), .C1(n3776), .Y(n431) );
  AOI222XL U4119 ( .A0(N798), .A1(n3782), .B0(N414), .B1(n250), .C0(N877), 
        .C1(n251), .Y(n432) );
  AND4X1 U4120 ( .A(n439), .B(n440), .C(n441), .D(n442), .Y(n143) );
  AOI221XL U4121 ( .A0(n443), .A1(n4015), .B0(n2677), .B1(n444), .C0(n445), 
        .Y(n442) );
  AOI222XL U4122 ( .A0(dataout[12]), .A1(n3772), .B0(N908), .B1(n253), .C0(
        N940), .C1(n3776), .Y(n439) );
  AOI222XL U4123 ( .A0(N797), .A1(n249), .B0(N413), .B1(n250), .C0(N876), .C1(
        n251), .Y(n440) );
  AND4X1 U4124 ( .A(n447), .B(n448), .C(n449), .D(n450), .Y(n144) );
  AOI221XL U4125 ( .A0(n451), .A1(n4016), .B0(n2676), .B1(n452), .C0(n453), 
        .Y(n450) );
  AOI222XL U4126 ( .A0(dataout[11]), .A1(n252), .B0(N907), .B1(n3777), .C0(
        N939), .C1(n3775), .Y(n447) );
  AOI222XL U4127 ( .A0(N796), .A1(n3782), .B0(N412), .B1(n3779), .C0(N875), 
        .C1(n3778), .Y(n448) );
  AND4X1 U4128 ( .A(n455), .B(n456), .C(n457), .D(n458), .Y(n145) );
  AOI221XL U4129 ( .A0(n459), .A1(n4017), .B0(n2673), .B1(n460), .C0(n461), 
        .Y(n458) );
  AOI222XL U4130 ( .A0(dataout[10]), .A1(n3771), .B0(N906), .B1(n253), .C0(
        N938), .C1(n3776), .Y(n455) );
  AOI222XL U4131 ( .A0(N795), .A1(n249), .B0(N411), .B1(n250), .C0(N874), .C1(
        n251), .Y(n456) );
  AND4X1 U4132 ( .A(n229), .B(n230), .C(n231), .D(n232), .Y(n113) );
  AOI221XL U4133 ( .A0(n233), .A1(n4018), .B0(n2674), .B1(n234), .C0(n235), 
        .Y(n232) );
  AOI222XL U4134 ( .A0(dataout[9]), .A1(n3772), .B0(N905), .B1(n253), .C0(N937), .C1(n3775), .Y(n229) );
  AOI222XL U4135 ( .A0(N794), .A1(n3782), .B0(N410), .B1(n250), .C0(N873), 
        .C1(n251), .Y(n230) );
  NOR2X1 U4136 ( .A(\R[3][22] ), .B(n3729), .Y(n3600) );
  NOR2X1 U4137 ( .A(\R[3][21] ), .B(n3729), .Y(n3605) );
  NOR2X1 U4138 ( .A(\R[3][20] ), .B(n3730), .Y(n3610) );
  NOR2X1 U4139 ( .A(\R[3][19] ), .B(n3730), .Y(n3615) );
  NOR2X1 U4140 ( .A(\R[3][18] ), .B(n3730), .Y(n3620) );
  NOR2X1 U4141 ( .A(n3747), .B(\R[1][22] ), .Y(n3602) );
  NOR2X1 U4142 ( .A(n3747), .B(\R[1][21] ), .Y(n3607) );
  NOR2X1 U4143 ( .A(n3747), .B(\R[1][20] ), .Y(n3612) );
  NOR2X1 U4144 ( .A(n3748), .B(\R[1][19] ), .Y(n3617) );
  NOR2X1 U4145 ( .A(n3748), .B(\R[1][18] ), .Y(n3622) );
  NOR2X1 U4146 ( .A(n3748), .B(\R[1][17] ), .Y(n3627) );
  AOI222XL U4147 ( .A0(dataout[3]), .A1(n3772), .B0(N899), .B1(n253), .C0(N931), .C1(n3775), .Y(n295) );
  MXI4X1 U4148 ( .A(\R[20][22] ), .B(\R[21][22] ), .C(\R[22][22] ), .D(
        \R[23][22] ), .S0(n3716), .S1(n3744), .Y(n3458) );
  MXI4X1 U4149 ( .A(\R[4][22] ), .B(\R[5][22] ), .C(\R[6][22] ), .D(\R[7][22] ), .S0(n3716), .S1(n3745), .Y(n3463) );
  MXI4X1 U4150 ( .A(\R[20][21] ), .B(\R[21][21] ), .C(\R[22][21] ), .D(
        \R[23][21] ), .S0(n3716), .S1(n3744), .Y(n3448) );
  MXI4X1 U4151 ( .A(\R[4][21] ), .B(\R[5][21] ), .C(\R[6][21] ), .D(\R[7][21] ), .S0(n3716), .S1(n3744), .Y(n3453) );
  MXI4X1 U4152 ( .A(\R[20][20] ), .B(\R[21][20] ), .C(\R[22][20] ), .D(
        \R[23][20] ), .S0(n3715), .S1(n3744), .Y(n3438) );
  MXI4X1 U4153 ( .A(\R[4][20] ), .B(\R[5][20] ), .C(\R[6][20] ), .D(\R[7][20] ), .S0(n3715), .S1(n3744), .Y(n3443) );
  MXI4X1 U4154 ( .A(\R[20][19] ), .B(\R[21][19] ), .C(\R[22][19] ), .D(
        \R[23][19] ), .S0(n3715), .S1(n3744), .Y(n3428) );
  MXI4X1 U4155 ( .A(\R[4][19] ), .B(\R[5][19] ), .C(\R[6][19] ), .D(\R[7][19] ), .S0(n3715), .S1(n3744), .Y(n3433) );
  MXI4X1 U4156 ( .A(\R[20][18] ), .B(\R[21][18] ), .C(\R[22][18] ), .D(
        \R[23][18] ), .S0(n3715), .S1(n3744), .Y(n3418) );
  MXI4X1 U4157 ( .A(\R[4][18] ), .B(\R[5][18] ), .C(\R[6][18] ), .D(\R[7][18] ), .S0(n3715), .S1(n3744), .Y(n3423) );
  MXI4X1 U4158 ( .A(\R[20][17] ), .B(\R[21][17] ), .C(\R[22][17] ), .D(
        \R[23][17] ), .S0(n3715), .S1(n3744), .Y(n3408) );
  MXI4X1 U4159 ( .A(\R[4][17] ), .B(\R[5][17] ), .C(\R[6][17] ), .D(\R[7][17] ), .S0(n3715), .S1(n3744), .Y(n3413) );
  MXI4X1 U4160 ( .A(\R[16][22] ), .B(\R[17][22] ), .C(\R[18][22] ), .D(
        \R[19][22] ), .S0(n3716), .S1(n3744), .Y(n3456) );
  MXI4X1 U4161 ( .A(\R[16][21] ), .B(\R[17][21] ), .C(\R[18][21] ), .D(
        \R[19][21] ), .S0(n3716), .S1(n3744), .Y(n3446) );
  MXI4X1 U4162 ( .A(\R[16][20] ), .B(\R[17][20] ), .C(\R[18][20] ), .D(
        \R[19][20] ), .S0(n3715), .S1(n3744), .Y(n3436) );
  MXI4X1 U4163 ( .A(\R[16][19] ), .B(\R[17][19] ), .C(\R[18][19] ), .D(
        \R[19][19] ), .S0(n3715), .S1(n3744), .Y(n3426) );
  MXI4X1 U4164 ( .A(\R[16][18] ), .B(\R[17][18] ), .C(\R[18][18] ), .D(
        \R[19][18] ), .S0(n3715), .S1(n3744), .Y(n3416) );
  MXI4X1 U4165 ( .A(\R[24][22] ), .B(\R[25][22] ), .C(\R[26][22] ), .D(
        \R[27][22] ), .S0(n3716), .S1(n3744), .Y(n3457) );
  MXI4X1 U4166 ( .A(\R[8][22] ), .B(\R[9][22] ), .C(\R[10][22] ), .D(
        \R[11][22] ), .S0(n3716), .S1(n3745), .Y(n3462) );
  MXI4X1 U4167 ( .A(\R[24][21] ), .B(\R[25][21] ), .C(\R[26][21] ), .D(
        \R[27][21] ), .S0(n3716), .S1(n3744), .Y(n3447) );
  MXI4X1 U4168 ( .A(\R[8][21] ), .B(\R[9][21] ), .C(\R[10][21] ), .D(
        \R[11][21] ), .S0(n3716), .S1(n3744), .Y(n3452) );
  MXI4X1 U4169 ( .A(\R[24][20] ), .B(\R[25][20] ), .C(\R[26][20] ), .D(
        \R[27][20] ), .S0(n3715), .S1(n3744), .Y(n3437) );
  MXI4X1 U4170 ( .A(\R[8][20] ), .B(\R[9][20] ), .C(\R[10][20] ), .D(
        \R[11][20] ), .S0(n3715), .S1(n3744), .Y(n3442) );
  MXI4X1 U4171 ( .A(\R[24][19] ), .B(\R[25][19] ), .C(\R[26][19] ), .D(
        \R[27][19] ), .S0(n3715), .S1(n3744), .Y(n3427) );
  MXI4X1 U4172 ( .A(\R[8][19] ), .B(\R[9][19] ), .C(\R[10][19] ), .D(
        \R[11][19] ), .S0(n3715), .S1(n3744), .Y(n3432) );
  MXI4X1 U4173 ( .A(\R[24][18] ), .B(\R[25][18] ), .C(\R[26][18] ), .D(
        \R[27][18] ), .S0(n3715), .S1(n3744), .Y(n3417) );
  MXI4X1 U4174 ( .A(\R[8][18] ), .B(\R[9][18] ), .C(\R[10][18] ), .D(
        \R[11][18] ), .S0(n3715), .S1(n3744), .Y(n3422) );
  MXI4X1 U4175 ( .A(\R[8][17] ), .B(\R[9][17] ), .C(\R[10][17] ), .D(
        \R[11][17] ), .S0(n3715), .S1(n3744), .Y(n3412) );
  MXI4X1 U4176 ( .A(\R[28][22] ), .B(\R[29][22] ), .C(\R[30][22] ), .D(
        \R[31][22] ), .S0(n3716), .S1(n3744), .Y(n3459) );
  MXI4X1 U4177 ( .A(\R[28][21] ), .B(\R[29][21] ), .C(\R[30][21] ), .D(
        \R[31][21] ), .S0(n3716), .S1(n3744), .Y(n3449) );
  MXI4X1 U4178 ( .A(\R[28][20] ), .B(\R[29][20] ), .C(\R[30][20] ), .D(
        \R[31][20] ), .S0(n3715), .S1(n3744), .Y(n3439) );
  MXI4X1 U4179 ( .A(\R[28][19] ), .B(\R[29][19] ), .C(\R[30][19] ), .D(
        \R[31][19] ), .S0(n3715), .S1(n3744), .Y(n3429) );
  MXI4X1 U4180 ( .A(\R[28][18] ), .B(\R[29][18] ), .C(\R[30][18] ), .D(
        \R[31][18] ), .S0(n3715), .S1(n3744), .Y(n3419) );
  MXI4X1 U4181 ( .A(\R[28][17] ), .B(\R[29][17] ), .C(\R[30][17] ), .D(
        \R[31][17] ), .S0(n3715), .S1(n3744), .Y(n3409) );
  OAI221XL U4182 ( .A0(n2728), .A1(n3783), .B0(n1574), .B1(n4045), .C0(n499), 
        .Y(n2608) );
  AOI22X1 U4183 ( .A0(N275), .A1(n3789), .B0(N1014), .B1(n3785), .Y(n499) );
  OAI221XL U4184 ( .A0(n4012), .A1(n478), .B0(n1575), .B1(n4045), .C0(n500), 
        .Y(n2609) );
  AOI22X1 U4185 ( .A0(N274), .A1(n3788), .B0(N1013), .B1(n3785), .Y(n500) );
  OAI221XL U4186 ( .A0(n4013), .A1(n478), .B0(n1576), .B1(n4045), .C0(n502), 
        .Y(n2610) );
  AOI22X1 U4187 ( .A0(N273), .A1(n3788), .B0(N1012), .B1(n3784), .Y(n502) );
  OAI221XL U4188 ( .A0(n2710), .A1(n3783), .B0(n1577), .B1(n4045), .C0(n503), 
        .Y(n2611) );
  AOI22X1 U4189 ( .A0(N272), .A1(n3788), .B0(N1011), .B1(n3784), .Y(n503) );
  OAI221XL U4190 ( .A0(n2716), .A1(n478), .B0(n1578), .B1(n4045), .C0(n504), 
        .Y(n2612) );
  AOI22X1 U4191 ( .A0(N271), .A1(n3788), .B0(N1010), .B1(n3784), .Y(n504) );
  OAI221XL U4192 ( .A0(n2713), .A1(n3783), .B0(n1579), .B1(n4045), .C0(n505), 
        .Y(n2613) );
  AOI22X1 U4193 ( .A0(N270), .A1(n3788), .B0(N1009), .B1(n3784), .Y(n505) );
  CLKMX2X2 U4194 ( .A(n3490), .B(n3485), .S0(n3769), .Y(N228) );
  MXI4X1 U4195 ( .A(n3491), .B(n3492), .C(n3493), .D(n3494), .S0(n3763), .S1(
        n3755), .Y(n3490) );
  MXI4X1 U4196 ( .A(n3486), .B(n3487), .C(n3488), .D(n3489), .S0(n3763), .S1(
        n3755), .Y(n3485) );
  MXI4X1 U4197 ( .A(\R[12][25] ), .B(\R[13][25] ), .C(\R[14][25] ), .D(
        \R[15][25] ), .S0(n3716), .S1(n3745), .Y(n3494) );
  CLKMX2X2 U4198 ( .A(n3470), .B(n3465), .S0(n3769), .Y(N230) );
  MXI4X1 U4199 ( .A(n3471), .B(n3472), .C(n3473), .D(n3474), .S0(n3763), .S1(
        n3755), .Y(n3470) );
  MXI4X1 U4200 ( .A(n3466), .B(n3467), .C(n3468), .D(n3469), .S0(n3763), .S1(
        n3755), .Y(n3465) );
  MXI4X1 U4201 ( .A(\R[12][23] ), .B(\R[13][23] ), .C(\R[14][23] ), .D(
        \R[15][23] ), .S0(n3716), .S1(n3745), .Y(n3474) );
  CLKMX2X2 U4202 ( .A(n3540), .B(n3535), .S0(n3769), .Y(N223) );
  MXI4X1 U4203 ( .A(n3541), .B(n3542), .C(n3543), .D(n3544), .S0(n3764), .S1(
        n3756), .Y(n3540) );
  MXI4X1 U4204 ( .A(n3536), .B(n3537), .C(n3538), .D(n3539), .S0(n3764), .S1(
        n3756), .Y(n3535) );
  MXI4X1 U4205 ( .A(\R[12][30] ), .B(\R[13][30] ), .C(\R[14][30] ), .D(
        \R[15][30] ), .S0(n3717), .S1(n3745), .Y(n3544) );
  CLKMX2X2 U4206 ( .A(n3500), .B(n3495), .S0(n3769), .Y(N227) );
  MXI4X1 U4207 ( .A(n3501), .B(n3502), .C(n3503), .D(n3504), .S0(n3764), .S1(
        n3756), .Y(n3500) );
  MXI4X1 U4208 ( .A(n3496), .B(n3497), .C(n3498), .D(n3499), .S0(n3764), .S1(
        n3756), .Y(n3495) );
  MXI4X1 U4209 ( .A(\R[12][26] ), .B(\R[13][26] ), .C(\R[14][26] ), .D(
        \R[15][26] ), .S0(n3716), .S1(n3745), .Y(n3504) );
  CLKMX2X2 U4210 ( .A(n3480), .B(n3475), .S0(n3769), .Y(N229) );
  MXI4X1 U4211 ( .A(n3481), .B(n3482), .C(n3483), .D(n3484), .S0(n3763), .S1(
        n3755), .Y(n3480) );
  MXI4X1 U4212 ( .A(n3476), .B(n3477), .C(n3478), .D(n3479), .S0(n3763), .S1(
        n3755), .Y(n3475) );
  MXI4X1 U4213 ( .A(\R[12][24] ), .B(\R[13][24] ), .C(\R[14][24] ), .D(
        \R[15][24] ), .S0(n3716), .S1(n3745), .Y(n3484) );
  CLKMX2X2 U4214 ( .A(n3520), .B(n3515), .S0(n3769), .Y(N225) );
  MXI4X1 U4215 ( .A(n3521), .B(n3522), .C(n3523), .D(n3524), .S0(n3764), .S1(
        n3756), .Y(n3520) );
  MXI4X1 U4216 ( .A(n3516), .B(n3517), .C(n3518), .D(n3519), .S0(n3764), .S1(
        n3756), .Y(n3515) );
  MXI4X1 U4217 ( .A(\R[12][28] ), .B(\R[13][28] ), .C(\R[14][28] ), .D(
        \R[15][28] ), .S0(n3716), .S1(n3745), .Y(n3524) );
  CLKMX2X2 U4218 ( .A(n3530), .B(n3525), .S0(n3769), .Y(N224) );
  MXI4X1 U4219 ( .A(n3531), .B(n3532), .C(n3533), .D(n3534), .S0(n3764), .S1(
        n3756), .Y(n3530) );
  MXI4X1 U4220 ( .A(n3526), .B(n3527), .C(n3528), .D(n3529), .S0(n3764), .S1(
        n3756), .Y(n3525) );
  MXI4X1 U4221 ( .A(\R[12][29] ), .B(\R[13][29] ), .C(\R[14][29] ), .D(
        \R[15][29] ), .S0(n3717), .S1(n3745), .Y(n3534) );
  CLKMX2X2 U4222 ( .A(n3550), .B(n3545), .S0(n3769), .Y(N222) );
  MXI4X1 U4223 ( .A(n3551), .B(n3552), .C(n3553), .D(n3554), .S0(n3764), .S1(
        n3756), .Y(n3550) );
  MXI4X1 U4224 ( .A(n3546), .B(n3547), .C(n3548), .D(n3549), .S0(n3764), .S1(
        n3756), .Y(n3545) );
  MXI4X1 U4225 ( .A(\R[12][31] ), .B(\R[13][31] ), .C(\R[14][31] ), .D(
        \R[15][31] ), .S0(n3717), .S1(n3745), .Y(n3554) );
  AOI222XL U4226 ( .A0(dataout[1]), .A1(n252), .B0(N897), .B1(n253), .C0(N929), 
        .C1(n3775), .Y(n385) );
  OAI22XL U4227 ( .A0(n3959), .A1(n168), .B0(n597), .B1(n3852), .Y(n1631) );
  OAI22XL U4228 ( .A0(n3956), .A1(n168), .B0(n598), .B1(n3852), .Y(n1632) );
  OAI22XL U4229 ( .A0(n3953), .A1(n168), .B0(n599), .B1(n3852), .Y(n1633) );
  OAI22XL U4230 ( .A0(n3950), .A1(n168), .B0(n600), .B1(n3852), .Y(n1634) );
  OAI22XL U4231 ( .A0(n3947), .A1(n168), .B0(n601), .B1(n3852), .Y(n1635) );
  OAI22XL U4232 ( .A0(n3935), .A1(n168), .B0(n603), .B1(n3852), .Y(n1637) );
  OAI22XL U4233 ( .A0(n3902), .A1(n168), .B0(n604), .B1(n3852), .Y(n1638) );
  OAI22XL U4234 ( .A0(n3870), .A1(n3851), .B0(n605), .B1(n3852), .Y(n1639) );
  OAI22XL U4235 ( .A0(n3959), .A1(n3849), .B0(n629), .B1(n3850), .Y(n1663) );
  OAI22XL U4236 ( .A0(n3956), .A1(n3849), .B0(n630), .B1(n3850), .Y(n1664) );
  OAI22XL U4237 ( .A0(n3953), .A1(n3849), .B0(n631), .B1(n3850), .Y(n1665) );
  OAI22XL U4238 ( .A0(n3950), .A1(n3849), .B0(n632), .B1(n3850), .Y(n1666) );
  OAI22XL U4239 ( .A0(n3947), .A1(n3849), .B0(n633), .B1(n3850), .Y(n1667) );
  OAI22XL U4240 ( .A0(n3935), .A1(n3849), .B0(n635), .B1(n3850), .Y(n1669) );
  OAI22XL U4241 ( .A0(n3902), .A1(n171), .B0(n636), .B1(n3850), .Y(n1670) );
  OAI22XL U4242 ( .A0(n3870), .A1(n171), .B0(n637), .B1(n3850), .Y(n1671) );
  OAI22XL U4243 ( .A0(n3959), .A1(n175), .B0(n661), .B1(n3845), .Y(n1695) );
  OAI22XL U4244 ( .A0(n3956), .A1(n175), .B0(n662), .B1(n3845), .Y(n1696) );
  OAI22XL U4245 ( .A0(n3953), .A1(n175), .B0(n663), .B1(n3845), .Y(n1697) );
  OAI22XL U4246 ( .A0(n3950), .A1(n175), .B0(n664), .B1(n3845), .Y(n1698) );
  OAI22XL U4247 ( .A0(n3947), .A1(n175), .B0(n665), .B1(n3845), .Y(n1699) );
  OAI22XL U4248 ( .A0(n3935), .A1(n175), .B0(n667), .B1(n3845), .Y(n1701) );
  OAI22XL U4249 ( .A0(n3902), .A1(n175), .B0(n668), .B1(n3845), .Y(n1702) );
  OAI22XL U4250 ( .A0(n3870), .A1(n3844), .B0(n669), .B1(n3845), .Y(n1703) );
  OAI22XL U4251 ( .A0(n3959), .A1(n3842), .B0(n693), .B1(n3843), .Y(n1727) );
  OAI22XL U4252 ( .A0(n3956), .A1(n3842), .B0(n694), .B1(n3843), .Y(n1728) );
  OAI22XL U4253 ( .A0(n3953), .A1(n3842), .B0(n695), .B1(n3843), .Y(n1729) );
  OAI22XL U4254 ( .A0(n3950), .A1(n3842), .B0(n696), .B1(n3843), .Y(n1730) );
  OAI22XL U4255 ( .A0(n3947), .A1(n3841), .B0(n697), .B1(n3843), .Y(n1731) );
  OAI22XL U4256 ( .A0(n3935), .A1(n3842), .B0(n699), .B1(n3843), .Y(n1733) );
  OAI22XL U4257 ( .A0(n3902), .A1(n177), .B0(n700), .B1(n3843), .Y(n1734) );
  OAI22XL U4258 ( .A0(n3870), .A1(n3841), .B0(n701), .B1(n3843), .Y(n1735) );
  OAI22XL U4259 ( .A0(n3960), .A1(n3839), .B0(n725), .B1(n3840), .Y(n1759) );
  OAI22XL U4260 ( .A0(n3957), .A1(n3839), .B0(n726), .B1(n3840), .Y(n1760) );
  OAI22XL U4261 ( .A0(n3954), .A1(n3839), .B0(n727), .B1(n3840), .Y(n1761) );
  OAI22XL U4262 ( .A0(n3951), .A1(n3839), .B0(n728), .B1(n3840), .Y(n1762) );
  OAI22XL U4263 ( .A0(n3948), .A1(n3839), .B0(n729), .B1(n3840), .Y(n1763) );
  OAI22XL U4264 ( .A0(n3936), .A1(n3839), .B0(n731), .B1(n3840), .Y(n1765) );
  OAI22XL U4265 ( .A0(n3903), .A1(n181), .B0(n732), .B1(n3840), .Y(n1766) );
  OAI22XL U4266 ( .A0(n3870), .A1(n181), .B0(n733), .B1(n3840), .Y(n1767) );
  OAI22XL U4267 ( .A0(n3960), .A1(n3837), .B0(n757), .B1(n3838), .Y(n1791) );
  OAI22XL U4268 ( .A0(n3957), .A1(n3837), .B0(n758), .B1(n3838), .Y(n1792) );
  OAI22XL U4269 ( .A0(n3954), .A1(n3837), .B0(n759), .B1(n3838), .Y(n1793) );
  OAI22XL U4270 ( .A0(n3951), .A1(n3837), .B0(n760), .B1(n3838), .Y(n1794) );
  OAI22XL U4271 ( .A0(n3948), .A1(n3837), .B0(n761), .B1(n3838), .Y(n1795) );
  OAI22XL U4272 ( .A0(n3936), .A1(n3837), .B0(n763), .B1(n3838), .Y(n1797) );
  OAI22XL U4273 ( .A0(n3903), .A1(n184), .B0(n764), .B1(n3838), .Y(n1798) );
  OAI22XL U4274 ( .A0(n3870), .A1(n184), .B0(n765), .B1(n3838), .Y(n1799) );
  OAI22XL U4275 ( .A0(n3960), .A1(n186), .B0(n789), .B1(n3836), .Y(n1823) );
  OAI22XL U4276 ( .A0(n3957), .A1(n186), .B0(n790), .B1(n3836), .Y(n1824) );
  OAI22XL U4277 ( .A0(n3954), .A1(n186), .B0(n791), .B1(n3836), .Y(n1825) );
  OAI22XL U4278 ( .A0(n3951), .A1(n186), .B0(n792), .B1(n3836), .Y(n1826) );
  OAI22XL U4279 ( .A0(n3948), .A1(n186), .B0(n793), .B1(n3836), .Y(n1827) );
  OAI22XL U4280 ( .A0(n3936), .A1(n186), .B0(n795), .B1(n3836), .Y(n1829) );
  OAI22XL U4281 ( .A0(n3903), .A1(n186), .B0(n796), .B1(n3836), .Y(n1830) );
  OAI22XL U4282 ( .A0(n3870), .A1(n3835), .B0(n797), .B1(n3836), .Y(n1831) );
  OAI22XL U4283 ( .A0(n3960), .A1(n3833), .B0(n821), .B1(n3834), .Y(n1855) );
  OAI22XL U4284 ( .A0(n3957), .A1(n3833), .B0(n822), .B1(n3834), .Y(n1856) );
  OAI22XL U4285 ( .A0(n3954), .A1(n3833), .B0(n823), .B1(n3834), .Y(n1857) );
  OAI22XL U4286 ( .A0(n3951), .A1(n3833), .B0(n824), .B1(n3834), .Y(n1858) );
  OAI22XL U4287 ( .A0(n3948), .A1(n3832), .B0(n825), .B1(n3834), .Y(n1859) );
  OAI22XL U4288 ( .A0(n3936), .A1(n3833), .B0(n827), .B1(n3834), .Y(n1861) );
  OAI22XL U4289 ( .A0(n3903), .A1(n188), .B0(n828), .B1(n3834), .Y(n1862) );
  OAI22XL U4290 ( .A0(n3870), .A1(n3832), .B0(n829), .B1(n3834), .Y(n1863) );
  OAI22XL U4291 ( .A0(n3960), .A1(n191), .B0(n853), .B1(n3831), .Y(n1887) );
  OAI22XL U4292 ( .A0(n3957), .A1(n191), .B0(n854), .B1(n3831), .Y(n1888) );
  OAI22XL U4293 ( .A0(n3954), .A1(n191), .B0(n855), .B1(n3831), .Y(n1889) );
  OAI22XL U4294 ( .A0(n3951), .A1(n191), .B0(n856), .B1(n3831), .Y(n1890) );
  OAI22XL U4295 ( .A0(n3948), .A1(n191), .B0(n857), .B1(n3831), .Y(n1891) );
  OAI22XL U4296 ( .A0(n3936), .A1(n191), .B0(n859), .B1(n3831), .Y(n1893) );
  OAI22XL U4297 ( .A0(n3903), .A1(n191), .B0(n860), .B1(n3831), .Y(n1894) );
  OAI22XL U4298 ( .A0(n3870), .A1(n3830), .B0(n861), .B1(n3831), .Y(n1895) );
  OAI22XL U4299 ( .A0(n3960), .A1(n3828), .B0(n885), .B1(n3829), .Y(n1919) );
  OAI22XL U4300 ( .A0(n3957), .A1(n3828), .B0(n886), .B1(n3829), .Y(n1920) );
  OAI22XL U4301 ( .A0(n3954), .A1(n3828), .B0(n887), .B1(n3829), .Y(n1921) );
  OAI22XL U4302 ( .A0(n3951), .A1(n3828), .B0(n888), .B1(n3829), .Y(n1922) );
  OAI22XL U4303 ( .A0(n3948), .A1(n3828), .B0(n889), .B1(n3829), .Y(n1923) );
  OAI22XL U4304 ( .A0(n3936), .A1(n3828), .B0(n891), .B1(n3829), .Y(n1925) );
  OAI22XL U4305 ( .A0(n3903), .A1(n194), .B0(n892), .B1(n3829), .Y(n1926) );
  OAI22XL U4306 ( .A0(n3870), .A1(n194), .B0(n893), .B1(n3829), .Y(n1927) );
  OAI22XL U4307 ( .A0(n3960), .A1(n196), .B0(n917), .B1(n3827), .Y(n1951) );
  OAI22XL U4308 ( .A0(n3957), .A1(n196), .B0(n918), .B1(n3827), .Y(n1952) );
  OAI22XL U4309 ( .A0(n3954), .A1(n196), .B0(n919), .B1(n3827), .Y(n1953) );
  OAI22XL U4310 ( .A0(n3951), .A1(n196), .B0(n920), .B1(n3827), .Y(n1954) );
  OAI22XL U4311 ( .A0(n3948), .A1(n196), .B0(n921), .B1(n3827), .Y(n1955) );
  OAI22XL U4312 ( .A0(n3936), .A1(n196), .B0(n923), .B1(n3827), .Y(n1957) );
  OAI22XL U4313 ( .A0(n3903), .A1(n196), .B0(n924), .B1(n3827), .Y(n1958) );
  OAI22XL U4314 ( .A0(n3870), .A1(n3826), .B0(n925), .B1(n3827), .Y(n1959) );
  OAI22XL U4315 ( .A0(n3960), .A1(n3824), .B0(n949), .B1(n3825), .Y(n1983) );
  OAI22XL U4316 ( .A0(n3957), .A1(n3824), .B0(n950), .B1(n3825), .Y(n1984) );
  OAI22XL U4317 ( .A0(n3954), .A1(n3824), .B0(n951), .B1(n3825), .Y(n1985) );
  OAI22XL U4318 ( .A0(n3951), .A1(n3824), .B0(n952), .B1(n3825), .Y(n1986) );
  OAI22XL U4319 ( .A0(n3948), .A1(n3823), .B0(n953), .B1(n3825), .Y(n1987) );
  OAI22XL U4320 ( .A0(n3936), .A1(n3824), .B0(n955), .B1(n3825), .Y(n1989) );
  OAI22XL U4321 ( .A0(n3903), .A1(n198), .B0(n956), .B1(n3825), .Y(n1990) );
  OAI22XL U4322 ( .A0(n3869), .A1(n3823), .B0(n957), .B1(n3825), .Y(n1991) );
  OAI22XL U4323 ( .A0(n3960), .A1(n204), .B0(n981), .B1(n3820), .Y(n2015) );
  OAI22XL U4324 ( .A0(n3957), .A1(n204), .B0(n982), .B1(n3820), .Y(n2016) );
  OAI22XL U4325 ( .A0(n3954), .A1(n204), .B0(n983), .B1(n3820), .Y(n2017) );
  OAI22XL U4326 ( .A0(n3951), .A1(n204), .B0(n984), .B1(n3820), .Y(n2018) );
  OAI22XL U4327 ( .A0(n3948), .A1(n204), .B0(n985), .B1(n3820), .Y(n2019) );
  OAI22XL U4328 ( .A0(n3936), .A1(n204), .B0(n987), .B1(n3820), .Y(n2021) );
  OAI22XL U4329 ( .A0(n3903), .A1(n204), .B0(n988), .B1(n3820), .Y(n2022) );
  OAI22XL U4330 ( .A0(n3869), .A1(n3819), .B0(n989), .B1(n3820), .Y(n2023) );
  OAI22XL U4331 ( .A0(n3960), .A1(n3817), .B0(n1013), .B1(n3818), .Y(n2047) );
  OAI22XL U4332 ( .A0(n3957), .A1(n3817), .B0(n1014), .B1(n3818), .Y(n2048) );
  OAI22XL U4333 ( .A0(n3954), .A1(n3817), .B0(n1015), .B1(n3818), .Y(n2049) );
  OAI22XL U4334 ( .A0(n3951), .A1(n3817), .B0(n1016), .B1(n3818), .Y(n2050) );
  OAI22XL U4335 ( .A0(n3948), .A1(n3817), .B0(n1017), .B1(n3818), .Y(n2051) );
  OAI22XL U4336 ( .A0(n3936), .A1(n3817), .B0(n1019), .B1(n3818), .Y(n2053) );
  OAI22XL U4337 ( .A0(n3903), .A1(n207), .B0(n1020), .B1(n3818), .Y(n2054) );
  OAI22XL U4338 ( .A0(n3869), .A1(n207), .B0(n1021), .B1(n3818), .Y(n2055) );
  OAI22XL U4339 ( .A0(n3960), .A1(n209), .B0(n1045), .B1(n3816), .Y(n2079) );
  OAI22XL U4340 ( .A0(n3957), .A1(n209), .B0(n1046), .B1(n3816), .Y(n2080) );
  OAI22XL U4341 ( .A0(n3954), .A1(n209), .B0(n1047), .B1(n3816), .Y(n2081) );
  OAI22XL U4342 ( .A0(n3951), .A1(n209), .B0(n1048), .B1(n3816), .Y(n2082) );
  OAI22XL U4343 ( .A0(n3948), .A1(n209), .B0(n1049), .B1(n3816), .Y(n2083) );
  OAI22XL U4344 ( .A0(n3936), .A1(n209), .B0(n1051), .B1(n3816), .Y(n2085) );
  OAI22XL U4345 ( .A0(n3903), .A1(n209), .B0(n1052), .B1(n3816), .Y(n2086) );
  OAI22XL U4346 ( .A0(n3869), .A1(n3815), .B0(n1053), .B1(n3816), .Y(n2087) );
  OAI22XL U4347 ( .A0(n3961), .A1(n3813), .B0(n1077), .B1(n3814), .Y(n2111) );
  OAI22XL U4348 ( .A0(n3958), .A1(n3813), .B0(n1078), .B1(n3814), .Y(n2112) );
  OAI22XL U4349 ( .A0(n3955), .A1(n3813), .B0(n1079), .B1(n3814), .Y(n2113) );
  OAI22XL U4350 ( .A0(n3952), .A1(n3813), .B0(n1080), .B1(n3814), .Y(n2114) );
  OAI22XL U4351 ( .A0(n3949), .A1(n3812), .B0(n1081), .B1(n3814), .Y(n2115) );
  OAI22XL U4352 ( .A0(n3937), .A1(n3813), .B0(n1083), .B1(n3814), .Y(n2117) );
  OAI22XL U4353 ( .A0(n3904), .A1(n211), .B0(n1084), .B1(n3814), .Y(n2118) );
  OAI22XL U4354 ( .A0(n3869), .A1(n3812), .B0(n1085), .B1(n3814), .Y(n2119) );
  OAI22XL U4355 ( .A0(n3961), .A1(n214), .B0(n1109), .B1(n3810), .Y(n2143) );
  OAI22XL U4356 ( .A0(n3958), .A1(n214), .B0(n1110), .B1(n3810), .Y(n2144) );
  OAI22XL U4357 ( .A0(n3955), .A1(n214), .B0(n1111), .B1(n3810), .Y(n2145) );
  OAI22XL U4358 ( .A0(n3952), .A1(n214), .B0(n1112), .B1(n3810), .Y(n2146) );
  OAI22XL U4359 ( .A0(n3949), .A1(n214), .B0(n1113), .B1(n3810), .Y(n2147) );
  OAI22XL U4360 ( .A0(n3937), .A1(n214), .B0(n1115), .B1(n3810), .Y(n2149) );
  OAI22XL U4361 ( .A0(n3904), .A1(n214), .B0(n1116), .B1(n3811), .Y(n2150) );
  OAI22XL U4362 ( .A0(n3869), .A1(n214), .B0(n1117), .B1(n3811), .Y(n2151) );
  OAI22XL U4363 ( .A0(n3961), .A1(n217), .B0(n1141), .B1(n3807), .Y(n2175) );
  OAI22XL U4364 ( .A0(n3958), .A1(n217), .B0(n1142), .B1(n3807), .Y(n2176) );
  OAI22XL U4365 ( .A0(n3955), .A1(n217), .B0(n1143), .B1(n3807), .Y(n2177) );
  OAI22XL U4366 ( .A0(n3952), .A1(n217), .B0(n1144), .B1(n3807), .Y(n2178) );
  OAI22XL U4367 ( .A0(n3949), .A1(n217), .B0(n1145), .B1(n3807), .Y(n2179) );
  OAI22XL U4368 ( .A0(n3937), .A1(n217), .B0(n1147), .B1(n3807), .Y(n2181) );
  OAI22XL U4369 ( .A0(n3904), .A1(n217), .B0(n1148), .B1(n3808), .Y(n2182) );
  OAI22XL U4370 ( .A0(n3869), .A1(n217), .B0(n1149), .B1(n3808), .Y(n2183) );
  OAI22XL U4371 ( .A0(n3961), .A1(n219), .B0(n1173), .B1(n3805), .Y(n2207) );
  OAI22XL U4372 ( .A0(n3958), .A1(n219), .B0(n1174), .B1(n3805), .Y(n2208) );
  OAI22XL U4373 ( .A0(n3955), .A1(n219), .B0(n1175), .B1(n3805), .Y(n2209) );
  OAI22XL U4374 ( .A0(n3952), .A1(n219), .B0(n1176), .B1(n3805), .Y(n2210) );
  OAI22XL U4375 ( .A0(n3949), .A1(n219), .B0(n1177), .B1(n3805), .Y(n2211) );
  OAI22XL U4376 ( .A0(n3937), .A1(n219), .B0(n1179), .B1(n3805), .Y(n2213) );
  OAI22XL U4377 ( .A0(n3904), .A1(n219), .B0(n1180), .B1(n3805), .Y(n2214) );
  OAI22XL U4378 ( .A0(n3869), .A1(n3804), .B0(n1181), .B1(n3805), .Y(n2215) );
  OAI22XL U4379 ( .A0(n3961), .A1(n222), .B0(n1205), .B1(n3802), .Y(n2239) );
  OAI22XL U4380 ( .A0(n3958), .A1(n222), .B0(n1206), .B1(n3802), .Y(n2240) );
  OAI22XL U4381 ( .A0(n3955), .A1(n222), .B0(n1207), .B1(n3802), .Y(n2241) );
  OAI22XL U4382 ( .A0(n3952), .A1(n222), .B0(n1208), .B1(n3802), .Y(n2242) );
  OAI22XL U4383 ( .A0(n3949), .A1(n222), .B0(n1209), .B1(n3802), .Y(n2243) );
  OAI22XL U4384 ( .A0(n3937), .A1(n222), .B0(n1211), .B1(n3802), .Y(n2245) );
  OAI22XL U4385 ( .A0(n3904), .A1(n222), .B0(n1212), .B1(n3803), .Y(n2246) );
  OAI22XL U4386 ( .A0(n3869), .A1(n222), .B0(n1213), .B1(n3803), .Y(n2247) );
  OAI22XL U4387 ( .A0(n3961), .A1(n225), .B0(n1237), .B1(n3800), .Y(n2271) );
  OAI22XL U4388 ( .A0(n3958), .A1(n225), .B0(n1238), .B1(n3800), .Y(n2272) );
  OAI22XL U4389 ( .A0(n3955), .A1(n225), .B0(n1239), .B1(n3800), .Y(n2273) );
  OAI22XL U4390 ( .A0(n3952), .A1(n225), .B0(n1240), .B1(n3800), .Y(n2274) );
  OAI22XL U4391 ( .A0(n3949), .A1(n225), .B0(n1241), .B1(n3800), .Y(n2275) );
  OAI22XL U4392 ( .A0(n3937), .A1(n225), .B0(n1243), .B1(n3800), .Y(n2277) );
  OAI22XL U4393 ( .A0(n3904), .A1(n225), .B0(n1244), .B1(n3800), .Y(n2278) );
  OAI22XL U4394 ( .A0(n3869), .A1(n3799), .B0(n1245), .B1(n3800), .Y(n2279) );
  OAI22XL U4395 ( .A0(n1269), .A1(n3798), .B0(n3961), .B1(n3795), .Y(n2303) );
  OAI22XL U4396 ( .A0(n1270), .A1(n3798), .B0(n3958), .B1(n3795), .Y(n2304) );
  OAI22XL U4397 ( .A0(n1271), .A1(n3798), .B0(n3955), .B1(n3795), .Y(n2305) );
  OAI22XL U4398 ( .A0(n1272), .A1(n3798), .B0(n3952), .B1(n3795), .Y(n2306) );
  OAI22XL U4399 ( .A0(n1273), .A1(n3798), .B0(n3949), .B1(n3796), .Y(n2307) );
  OAI22XL U4400 ( .A0(n1275), .A1(n3798), .B0(n3937), .B1(n3796), .Y(n2309) );
  OAI22XL U4401 ( .A0(n1276), .A1(n3798), .B0(n3904), .B1(n3797), .Y(n2310) );
  OAI22XL U4402 ( .A0(n3869), .A1(n3794), .B0(n1277), .B1(n3798), .Y(n2311) );
  OAI22XL U4403 ( .A0(n3959), .A1(n114), .B0(n1301), .B1(n3963), .Y(n2335) );
  OAI22XL U4404 ( .A0(n3956), .A1(n114), .B0(n1302), .B1(n3963), .Y(n2336) );
  OAI22XL U4405 ( .A0(n3953), .A1(n114), .B0(n1303), .B1(n3963), .Y(n2337) );
  OAI22XL U4406 ( .A0(n3950), .A1(n114), .B0(n1304), .B1(n3963), .Y(n2338) );
  OAI22XL U4407 ( .A0(n3947), .A1(n114), .B0(n1305), .B1(n3963), .Y(n2339) );
  OAI22XL U4408 ( .A0(n3935), .A1(n114), .B0(n1307), .B1(n3963), .Y(n2341) );
  OAI22XL U4409 ( .A0(n3902), .A1(n114), .B0(n1308), .B1(n3963), .Y(n2342) );
  OAI22XL U4410 ( .A0(n3871), .A1(n3962), .B0(n1309), .B1(n3963), .Y(n2343) );
  OAI22XL U4411 ( .A0(n3959), .A1(n149), .B0(n1333), .B1(n3868), .Y(n2367) );
  OAI22XL U4412 ( .A0(n3956), .A1(n149), .B0(n1334), .B1(n3868), .Y(n2368) );
  OAI22XL U4413 ( .A0(n3953), .A1(n149), .B0(n1335), .B1(n3868), .Y(n2369) );
  OAI22XL U4414 ( .A0(n3950), .A1(n149), .B0(n1336), .B1(n3868), .Y(n2370) );
  OAI22XL U4415 ( .A0(n3947), .A1(n149), .B0(n1337), .B1(n3868), .Y(n2371) );
  OAI22XL U4416 ( .A0(n3935), .A1(n149), .B0(n1339), .B1(n3868), .Y(n2373) );
  OAI22XL U4417 ( .A0(n3902), .A1(n149), .B0(n1340), .B1(n3868), .Y(n2374) );
  OAI22XL U4418 ( .A0(n3871), .A1(n3867), .B0(n1341), .B1(n3868), .Y(n2375) );
  OAI22XL U4419 ( .A0(n3959), .A1(n152), .B0(n1365), .B1(n3865), .Y(n2399) );
  OAI22XL U4420 ( .A0(n3956), .A1(n152), .B0(n1366), .B1(n3865), .Y(n2400) );
  OAI22XL U4421 ( .A0(n3953), .A1(n152), .B0(n1367), .B1(n3865), .Y(n2401) );
  OAI22XL U4422 ( .A0(n3950), .A1(n152), .B0(n1368), .B1(n3865), .Y(n2402) );
  OAI22XL U4423 ( .A0(n3947), .A1(n152), .B0(n1369), .B1(n3865), .Y(n2403) );
  OAI22XL U4424 ( .A0(n3935), .A1(n152), .B0(n1371), .B1(n3865), .Y(n2405) );
  OAI22XL U4425 ( .A0(n3902), .A1(n152), .B0(n1372), .B1(n3866), .Y(n2406) );
  OAI22XL U4426 ( .A0(n3871), .A1(n152), .B0(n1373), .B1(n3866), .Y(n2407) );
  OAI22XL U4427 ( .A0(n3959), .A1(n156), .B0(n1397), .B1(n3862), .Y(n2431) );
  OAI22XL U4428 ( .A0(n3956), .A1(n156), .B0(n1398), .B1(n3862), .Y(n2432) );
  OAI22XL U4429 ( .A0(n3953), .A1(n156), .B0(n1399), .B1(n3862), .Y(n2433) );
  OAI22XL U4430 ( .A0(n3950), .A1(n156), .B0(n1400), .B1(n3862), .Y(n2434) );
  OAI22XL U4431 ( .A0(n3947), .A1(n156), .B0(n1401), .B1(n3862), .Y(n2435) );
  OAI22XL U4432 ( .A0(n3935), .A1(n156), .B0(n1403), .B1(n3862), .Y(n2437) );
  OAI22XL U4433 ( .A0(n3902), .A1(n156), .B0(n1404), .B1(n3863), .Y(n2438) );
  OAI22XL U4434 ( .A0(n3871), .A1(n156), .B0(n1405), .B1(n3863), .Y(n2439) );
  OAI22XL U4435 ( .A0(n3959), .A1(n159), .B0(n1429), .B1(n3859), .Y(n2463) );
  OAI22XL U4436 ( .A0(n3956), .A1(n159), .B0(n1430), .B1(n3859), .Y(n2464) );
  OAI22XL U4437 ( .A0(n3953), .A1(n159), .B0(n1431), .B1(n3859), .Y(n2465) );
  OAI22XL U4438 ( .A0(n3950), .A1(n159), .B0(n1432), .B1(n3859), .Y(n2466) );
  OAI22XL U4439 ( .A0(n3947), .A1(n159), .B0(n1433), .B1(n3859), .Y(n2467) );
  OAI22XL U4440 ( .A0(n3935), .A1(n159), .B0(n1435), .B1(n3859), .Y(n2469) );
  OAI22XL U4441 ( .A0(n3902), .A1(n159), .B0(n1436), .B1(n3860), .Y(n2470) );
  OAI22XL U4442 ( .A0(n3871), .A1(n159), .B0(n1437), .B1(n3860), .Y(n2471) );
  OAI22XL U4443 ( .A0(n3959), .A1(n161), .B0(n1461), .B1(n3856), .Y(n2495) );
  OAI22XL U4444 ( .A0(n3956), .A1(n161), .B0(n1462), .B1(n3856), .Y(n2496) );
  OAI22XL U4445 ( .A0(n3953), .A1(n161), .B0(n1463), .B1(n3856), .Y(n2497) );
  OAI22XL U4446 ( .A0(n3950), .A1(n161), .B0(n1464), .B1(n3856), .Y(n2498) );
  OAI22XL U4447 ( .A0(n3947), .A1(n161), .B0(n1465), .B1(n3856), .Y(n2499) );
  OAI22XL U4448 ( .A0(n3935), .A1(n161), .B0(n1467), .B1(n3856), .Y(n2501) );
  OAI22XL U4449 ( .A0(n3902), .A1(n161), .B0(n1468), .B1(n3857), .Y(n2502) );
  OAI22XL U4450 ( .A0(n3871), .A1(n161), .B0(n1469), .B1(n3857), .Y(n2503) );
  OAI22XL U4451 ( .A0(n3959), .A1(n165), .B0(n1493), .B1(n3854), .Y(n2527) );
  OAI22XL U4452 ( .A0(n3956), .A1(n165), .B0(n1494), .B1(n3854), .Y(n2528) );
  OAI22XL U4453 ( .A0(n3953), .A1(n165), .B0(n1495), .B1(n3854), .Y(n2529) );
  OAI22XL U4454 ( .A0(n3950), .A1(n165), .B0(n1496), .B1(n3854), .Y(n2530) );
  OAI22XL U4455 ( .A0(n3947), .A1(n165), .B0(n1497), .B1(n3854), .Y(n2531) );
  OAI22XL U4456 ( .A0(n3935), .A1(n165), .B0(n1499), .B1(n3854), .Y(n2533) );
  OAI22XL U4457 ( .A0(n3902), .A1(n165), .B0(n1500), .B1(n3854), .Y(n2534) );
  OAI22XL U4458 ( .A0(n3871), .A1(n3853), .B0(n1501), .B1(n3854), .Y(n2535) );
  OAI22XL U4459 ( .A0(n3959), .A1(n3847), .B0(n1525), .B1(n3848), .Y(n2559) );
  OAI22XL U4460 ( .A0(n3956), .A1(n3847), .B0(n1526), .B1(n3848), .Y(n2560) );
  OAI22XL U4461 ( .A0(n3953), .A1(n3847), .B0(n1527), .B1(n3848), .Y(n2561) );
  OAI22XL U4462 ( .A0(n3950), .A1(n3847), .B0(n1528), .B1(n3848), .Y(n2562) );
  OAI22XL U4463 ( .A0(n3947), .A1(n3847), .B0(n1529), .B1(n3848), .Y(n2563) );
  OAI22XL U4464 ( .A0(n3935), .A1(n3846), .B0(n1531), .B1(n3848), .Y(n2565) );
  OAI22XL U4465 ( .A0(n3902), .A1(n173), .B0(n1532), .B1(n3848), .Y(n2566) );
  OAI22XL U4466 ( .A0(n3870), .A1(n3846), .B0(n1533), .B1(n3848), .Y(n2567) );
  OAI22XL U4467 ( .A0(n3960), .A1(n201), .B0(n1557), .B1(n3822), .Y(n2591) );
  OAI22XL U4468 ( .A0(n3957), .A1(n201), .B0(n1558), .B1(n3822), .Y(n2592) );
  OAI22XL U4469 ( .A0(n3954), .A1(n201), .B0(n1559), .B1(n3822), .Y(n2593) );
  OAI22XL U4470 ( .A0(n3951), .A1(n201), .B0(n1560), .B1(n3822), .Y(n2594) );
  OAI22XL U4471 ( .A0(n3948), .A1(n201), .B0(n1561), .B1(n3822), .Y(n2595) );
  OAI22XL U4472 ( .A0(n3936), .A1(n201), .B0(n1563), .B1(n3822), .Y(n2597) );
  OAI22XL U4473 ( .A0(n3903), .A1(n201), .B0(n1564), .B1(n3822), .Y(n2598) );
  OAI22XL U4474 ( .A0(n3869), .A1(n3821), .B0(n1565), .B1(n3822), .Y(n2599) );
  AND4X1 U4475 ( .A(n255), .B(n256), .C(n257), .D(n258), .Y(n116) );
  AOI221XL U4476 ( .A0(n259), .A1(n4019), .B0(n2675), .B1(n260), .C0(n261), 
        .Y(n258) );
  AOI222XL U4477 ( .A0(dataout[8]), .A1(n3772), .B0(N904), .B1(n253), .C0(N936), .C1(n3776), .Y(n255) );
  AOI222XL U4478 ( .A0(N793), .A1(n249), .B0(N409), .B1(n250), .C0(N872), .C1(
        n251), .Y(n256) );
  AND4X1 U4479 ( .A(n263), .B(n264), .C(n265), .D(n266), .Y(n117) );
  AOI221XL U4480 ( .A0(n267), .A1(n4020), .B0(n2671), .B1(n268), .C0(n269), 
        .Y(n266) );
  AOI222XL U4481 ( .A0(dataout[7]), .A1(n252), .B0(N903), .B1(n253), .C0(N935), 
        .C1(n3775), .Y(n263) );
  AOI222XL U4482 ( .A0(N792), .A1(n3782), .B0(N408), .B1(n250), .C0(N871), 
        .C1(n251), .Y(n264) );
  AND4X1 U4483 ( .A(n271), .B(n272), .C(n273), .D(n274), .Y(n118) );
  AOI221XL U4484 ( .A0(n275), .A1(n4021), .B0(n2672), .B1(n276), .C0(n277), 
        .Y(n274) );
  AOI222XL U4485 ( .A0(dataout[6]), .A1(n3772), .B0(N902), .B1(n253), .C0(N934), .C1(n3775), .Y(n271) );
  AOI222XL U4486 ( .A0(N791), .A1(n249), .B0(N407), .B1(n250), .C0(N870), .C1(
        n251), .Y(n272) );
  AND4X1 U4487 ( .A(n279), .B(n280), .C(n281), .D(n282), .Y(n119) );
  AOI221XL U4488 ( .A0(n283), .A1(n4022), .B0(n2655), .B1(n284), .C0(n285), 
        .Y(n282) );
  AOI222XL U4489 ( .A0(dataout[5]), .A1(n3772), .B0(N901), .B1(n253), .C0(N933), .C1(n3776), .Y(n279) );
  AOI222XL U4490 ( .A0(N790), .A1(n3782), .B0(N406), .B1(n250), .C0(N869), 
        .C1(n251), .Y(n280) );
  AND4X1 U4491 ( .A(n466), .B(n467), .C(n468), .D(n469), .Y(n146) );
  AOI222XL U4492 ( .A0(N593), .A1(n248), .B0(N253), .B1(n462), .C0(N657), .C1(
        n247), .Y(n468) );
  AOI221XL U4493 ( .A0(N864), .A1(n251), .B0(N785), .B1(n249), .C0(n477), .Y(
        n467) );
  AOI222XL U4494 ( .A0(dataout[0]), .A1(n3772), .B0(N896), .B1(n3777), .C0(
        N928), .C1(n3775), .Y(n466) );
  NOR2X1 U4495 ( .A(\R[3][31] ), .B(n3727), .Y(n3555) );
  NOR2X1 U4496 ( .A(\R[3][30] ), .B(n3727), .Y(n3560) );
  NOR2X1 U4497 ( .A(\R[3][29] ), .B(n3727), .Y(n3565) );
  NOR2X1 U4498 ( .A(\R[3][28] ), .B(n3728), .Y(n3570) );
  NOR2X1 U4499 ( .A(\R[3][27] ), .B(n3728), .Y(n3575) );
  NOR2X1 U4500 ( .A(\R[3][26] ), .B(n3728), .Y(n3580) );
  NOR2X1 U4501 ( .A(\R[3][25] ), .B(n3728), .Y(n3585) );
  NOR2X1 U4502 ( .A(\R[3][24] ), .B(n3729), .Y(n3590) );
  NOR2X1 U4503 ( .A(\R[3][23] ), .B(n3729), .Y(n3595) );
  NOR2X1 U4504 ( .A(n3747), .B(\R[1][25] ), .Y(n3587) );
  NOR2X1 U4505 ( .A(n3747), .B(\R[1][24] ), .Y(n3592) );
  NOR2X1 U4506 ( .A(n3747), .B(\R[1][23] ), .Y(n3597) );
  NOR2X1 U4507 ( .A(n3746), .B(\R[1][31] ), .Y(n3557) );
  NOR2X1 U4508 ( .A(n3746), .B(\R[1][30] ), .Y(n3562) );
  NOR2X1 U4509 ( .A(n3746), .B(\R[1][29] ), .Y(n3567) );
  NOR2X1 U4510 ( .A(n3746), .B(\R[1][28] ), .Y(n3572) );
  NOR2X1 U4511 ( .A(n3746), .B(\R[1][27] ), .Y(n3577) );
  NOR2X1 U4512 ( .A(n3746), .B(\R[1][26] ), .Y(n3582) );
  CLKMX2X2 U4513 ( .A(n3510), .B(n3505), .S0(n3769), .Y(N226) );
  MXI4X1 U4514 ( .A(n3511), .B(n3512), .C(n3513), .D(n3514), .S0(n3764), .S1(
        n3756), .Y(n3510) );
  MXI4X1 U4515 ( .A(n3506), .B(n3507), .C(n3508), .D(n3509), .S0(n3764), .S1(
        n3756), .Y(n3505) );
  MXI4X1 U4516 ( .A(\R[12][27] ), .B(\R[13][27] ), .C(\R[14][27] ), .D(
        \R[15][27] ), .S0(n3716), .S1(n3745), .Y(n3514) );
  AOI222XL U4517 ( .A0(dataout[2]), .A1(n3772), .B0(N898), .B1(n253), .C0(N930), .C1(n3776), .Y(n317) );
  AOI222XL U4518 ( .A0(dataout[4]), .A1(n252), .B0(N900), .B1(n253), .C0(N932), 
        .C1(n3776), .Y(n287) );
  MXI4X1 U4519 ( .A(\R[20][31] ), .B(\R[21][31] ), .C(\R[22][31] ), .D(
        \R[23][31] ), .S0(n3717), .S1(n3745), .Y(n3548) );
  MXI4X1 U4520 ( .A(\R[4][31] ), .B(\R[5][31] ), .C(\R[6][31] ), .D(\R[7][31] ), .S0(n3719), .S1(n3746), .Y(n3553) );
  MXI4X1 U4521 ( .A(\R[20][30] ), .B(\R[21][30] ), .C(\R[22][30] ), .D(
        \R[23][30] ), .S0(n3717), .S1(n3745), .Y(n3538) );
  MXI4X1 U4522 ( .A(\R[4][30] ), .B(\R[5][30] ), .C(\R[6][30] ), .D(\R[7][30] ), .S0(n3717), .S1(n3745), .Y(n3543) );
  MXI4X1 U4523 ( .A(\R[20][29] ), .B(\R[21][29] ), .C(\R[22][29] ), .D(
        \R[23][29] ), .S0(n3717), .S1(n3745), .Y(n3528) );
  MXI4X1 U4524 ( .A(\R[4][29] ), .B(\R[5][29] ), .C(\R[6][29] ), .D(\R[7][29] ), .S0(n3717), .S1(n3745), .Y(n3533) );
  MXI4X1 U4525 ( .A(\R[20][28] ), .B(\R[21][28] ), .C(\R[22][28] ), .D(
        \R[23][28] ), .S0(n3716), .S1(n3745), .Y(n3518) );
  MXI4X1 U4526 ( .A(\R[4][28] ), .B(\R[5][28] ), .C(\R[6][28] ), .D(\R[7][28] ), .S0(n3716), .S1(n3745), .Y(n3523) );
  MXI4X1 U4527 ( .A(\R[20][27] ), .B(\R[21][27] ), .C(\R[22][27] ), .D(
        \R[23][27] ), .S0(n3716), .S1(n3745), .Y(n3508) );
  MXI4X1 U4528 ( .A(\R[4][27] ), .B(\R[5][27] ), .C(\R[6][27] ), .D(\R[7][27] ), .S0(n3716), .S1(n3745), .Y(n3513) );
  MXI4X1 U4529 ( .A(\R[20][26] ), .B(\R[21][26] ), .C(\R[22][26] ), .D(
        \R[23][26] ), .S0(n3716), .S1(n3745), .Y(n3498) );
  MXI4X1 U4530 ( .A(\R[4][26] ), .B(\R[5][26] ), .C(\R[6][26] ), .D(\R[7][26] ), .S0(n3716), .S1(n3745), .Y(n3503) );
  MXI4X1 U4531 ( .A(\R[20][25] ), .B(\R[21][25] ), .C(\R[22][25] ), .D(
        \R[23][25] ), .S0(n3716), .S1(n3745), .Y(n3488) );
  MXI4X1 U4532 ( .A(\R[4][25] ), .B(\R[5][25] ), .C(\R[6][25] ), .D(\R[7][25] ), .S0(n3716), .S1(n3745), .Y(n3493) );
  MXI4X1 U4533 ( .A(\R[20][24] ), .B(\R[21][24] ), .C(\R[22][24] ), .D(
        \R[23][24] ), .S0(n3716), .S1(n3745), .Y(n3478) );
  MXI4X1 U4534 ( .A(\R[4][24] ), .B(\R[5][24] ), .C(\R[6][24] ), .D(\R[7][24] ), .S0(n3716), .S1(n3745), .Y(n3483) );
  MXI4X1 U4535 ( .A(\R[20][23] ), .B(\R[21][23] ), .C(\R[22][23] ), .D(
        \R[23][23] ), .S0(n3716), .S1(n3745), .Y(n3468) );
  MXI4X1 U4536 ( .A(\R[4][23] ), .B(\R[5][23] ), .C(\R[6][23] ), .D(\R[7][23] ), .S0(n3716), .S1(n3745), .Y(n3473) );
  MXI4X1 U4537 ( .A(\R[16][31] ), .B(\R[17][31] ), .C(\R[18][31] ), .D(
        \R[19][31] ), .S0(n3717), .S1(n3745), .Y(n3546) );
  MXI4X1 U4538 ( .A(\R[16][30] ), .B(\R[17][30] ), .C(\R[18][30] ), .D(
        \R[19][30] ), .S0(n3717), .S1(n3745), .Y(n3536) );
  MXI4X1 U4539 ( .A(\R[16][29] ), .B(\R[17][29] ), .C(\R[18][29] ), .D(
        \R[19][29] ), .S0(n3717), .S1(n3745), .Y(n3526) );
  MXI4X1 U4540 ( .A(\R[16][28] ), .B(\R[17][28] ), .C(\R[18][28] ), .D(
        \R[19][28] ), .S0(n3716), .S1(n3745), .Y(n3516) );
  MXI4X1 U4541 ( .A(\R[16][27] ), .B(\R[17][27] ), .C(\R[18][27] ), .D(
        \R[19][27] ), .S0(n3716), .S1(n3745), .Y(n3506) );
  MXI4X1 U4542 ( .A(\R[16][26] ), .B(\R[17][26] ), .C(\R[18][26] ), .D(
        \R[19][26] ), .S0(n3716), .S1(n3745), .Y(n3496) );
  MXI4X1 U4543 ( .A(\R[16][25] ), .B(\R[17][25] ), .C(\R[18][25] ), .D(
        \R[19][25] ), .S0(n3716), .S1(n3745), .Y(n3486) );
  MXI4X1 U4544 ( .A(\R[16][24] ), .B(\R[17][24] ), .C(\R[18][24] ), .D(
        \R[19][24] ), .S0(n3716), .S1(n3745), .Y(n3476) );
  MXI4X1 U4545 ( .A(\R[16][23] ), .B(\R[17][23] ), .C(\R[18][23] ), .D(
        \R[19][23] ), .S0(n3716), .S1(n3745), .Y(n3466) );
  MXI4X1 U4546 ( .A(\R[24][31] ), .B(\R[25][31] ), .C(\R[26][31] ), .D(
        \R[27][31] ), .S0(n3717), .S1(n3745), .Y(n3547) );
  MXI4X1 U4547 ( .A(\R[8][31] ), .B(\R[9][31] ), .C(\R[10][31] ), .D(
        \R[11][31] ), .S0(n3716), .S1(n3745), .Y(n3552) );
  MXI4X1 U4548 ( .A(\R[24][30] ), .B(\R[25][30] ), .C(\R[26][30] ), .D(
        \R[27][30] ), .S0(n3717), .S1(n3745), .Y(n3537) );
  MXI4X1 U4549 ( .A(\R[8][30] ), .B(\R[9][30] ), .C(\R[10][30] ), .D(
        \R[11][30] ), .S0(n3717), .S1(n3745), .Y(n3542) );
  MXI4X1 U4550 ( .A(\R[24][29] ), .B(\R[25][29] ), .C(\R[26][29] ), .D(
        \R[27][29] ), .S0(n3717), .S1(n3745), .Y(n3527) );
  MXI4X1 U4551 ( .A(\R[8][29] ), .B(\R[9][29] ), .C(\R[10][29] ), .D(
        \R[11][29] ), .S0(n3717), .S1(n3745), .Y(n3532) );
  MXI4X1 U4552 ( .A(\R[24][28] ), .B(\R[25][28] ), .C(\R[26][28] ), .D(
        \R[27][28] ), .S0(n3716), .S1(n3745), .Y(n3517) );
  MXI4X1 U4553 ( .A(\R[8][28] ), .B(\R[9][28] ), .C(\R[10][28] ), .D(
        \R[11][28] ), .S0(n3716), .S1(n3745), .Y(n3522) );
  MXI4X1 U4554 ( .A(\R[24][27] ), .B(\R[25][27] ), .C(\R[26][27] ), .D(
        \R[27][27] ), .S0(n3716), .S1(n3745), .Y(n3507) );
  MXI4X1 U4555 ( .A(\R[8][27] ), .B(\R[9][27] ), .C(\R[10][27] ), .D(
        \R[11][27] ), .S0(n3716), .S1(n3745), .Y(n3512) );
  MXI4X1 U4556 ( .A(\R[24][26] ), .B(\R[25][26] ), .C(\R[26][26] ), .D(
        \R[27][26] ), .S0(n3716), .S1(n3745), .Y(n3497) );
  MXI4X1 U4557 ( .A(\R[8][26] ), .B(\R[9][26] ), .C(\R[10][26] ), .D(
        \R[11][26] ), .S0(n3716), .S1(n3745), .Y(n3502) );
  MXI4X1 U4558 ( .A(\R[24][25] ), .B(\R[25][25] ), .C(\R[26][25] ), .D(
        \R[27][25] ), .S0(n3716), .S1(n3745), .Y(n3487) );
  MXI4X1 U4559 ( .A(\R[8][25] ), .B(\R[9][25] ), .C(\R[10][25] ), .D(
        \R[11][25] ), .S0(n3716), .S1(n3745), .Y(n3492) );
  MXI4X1 U4560 ( .A(\R[24][24] ), .B(\R[25][24] ), .C(\R[26][24] ), .D(
        \R[27][24] ), .S0(n3716), .S1(n3745), .Y(n3477) );
  MXI4X1 U4561 ( .A(\R[8][24] ), .B(\R[9][24] ), .C(\R[10][24] ), .D(
        \R[11][24] ), .S0(n3716), .S1(n3745), .Y(n3482) );
  MXI4X1 U4562 ( .A(\R[24][23] ), .B(\R[25][23] ), .C(\R[26][23] ), .D(
        \R[27][23] ), .S0(n3716), .S1(n3745), .Y(n3467) );
  MXI4X1 U4563 ( .A(\R[8][23] ), .B(\R[9][23] ), .C(\R[10][23] ), .D(
        \R[11][23] ), .S0(n3716), .S1(n3745), .Y(n3472) );
  MXI4X1 U4564 ( .A(\R[28][31] ), .B(\R[29][31] ), .C(\R[30][31] ), .D(
        \R[31][31] ), .S0(n3717), .S1(n3745), .Y(n3549) );
  MXI4X1 U4565 ( .A(\R[28][30] ), .B(\R[29][30] ), .C(\R[30][30] ), .D(
        \R[31][30] ), .S0(n3717), .S1(n3745), .Y(n3539) );
  MXI4X1 U4566 ( .A(\R[28][29] ), .B(\R[29][29] ), .C(\R[30][29] ), .D(
        \R[31][29] ), .S0(n3716), .S1(n3745), .Y(n3529) );
  MXI4X1 U4567 ( .A(\R[28][28] ), .B(\R[29][28] ), .C(\R[30][28] ), .D(
        \R[31][28] ), .S0(n3716), .S1(n3745), .Y(n3519) );
  MXI4X1 U4568 ( .A(\R[28][27] ), .B(\R[29][27] ), .C(\R[30][27] ), .D(
        \R[31][27] ), .S0(n3716), .S1(n3745), .Y(n3509) );
  MXI4X1 U4569 ( .A(\R[28][26] ), .B(\R[29][26] ), .C(\R[30][26] ), .D(
        \R[31][26] ), .S0(n3716), .S1(n3745), .Y(n3499) );
  MXI4X1 U4570 ( .A(\R[28][25] ), .B(\R[29][25] ), .C(\R[30][25] ), .D(
        \R[31][25] ), .S0(n3716), .S1(n3745), .Y(n3489) );
  MXI4X1 U4571 ( .A(\R[28][24] ), .B(\R[29][24] ), .C(\R[30][24] ), .D(
        \R[31][24] ), .S0(n3716), .S1(n3745), .Y(n3479) );
  MXI4X1 U4572 ( .A(\R[28][23] ), .B(\R[29][23] ), .C(\R[30][23] ), .D(
        \R[31][23] ), .S0(n3716), .S1(n3745), .Y(n3469) );
  OAI221XL U4573 ( .A0(n4014), .A1(n478), .B0(n1580), .B1(n4045), .C0(n506), 
        .Y(n2614) );
  AOI22X1 U4574 ( .A0(N269), .A1(n3788), .B0(N1008), .B1(n3784), .Y(n506) );
  OAI221XL U4575 ( .A0(n2750), .A1(n3783), .B0(n1581), .B1(n4045), .C0(n507), 
        .Y(n2615) );
  AOI22X1 U4576 ( .A0(N268), .A1(n3788), .B0(N1007), .B1(n3784), .Y(n507) );
  OAI221XL U4577 ( .A0(n2741), .A1(n478), .B0(n1582), .B1(n4045), .C0(n508), 
        .Y(n2616) );
  AOI22X1 U4578 ( .A0(N267), .A1(n3788), .B0(N1006), .B1(n3784), .Y(n508) );
  OAI221XL U4579 ( .A0(n4015), .A1(n3783), .B0(n1583), .B1(n4045), .C0(n509), 
        .Y(n2617) );
  AOI22X1 U4580 ( .A0(N266), .A1(n3788), .B0(N1005), .B1(n3784), .Y(n509) );
  OAI221XL U4581 ( .A0(n4016), .A1(n478), .B0(n1584), .B1(n4045), .C0(n510), 
        .Y(n2618) );
  AOI22X1 U4582 ( .A0(N265), .A1(n3788), .B0(N1004), .B1(n3784), .Y(n510) );
  OAI221XL U4583 ( .A0(n4017), .A1(n3783), .B0(n1585), .B1(n4045), .C0(n511), 
        .Y(n2619) );
  AOI22X1 U4584 ( .A0(N264), .A1(n3788), .B0(N1003), .B1(n3784), .Y(n511) );
  OAI221XL U4585 ( .A0(n4018), .A1(n3783), .B0(n1586), .B1(n4045), .C0(n479), 
        .Y(n2620) );
  AOI22X1 U4586 ( .A0(N263), .A1(n3790), .B0(N1002), .B1(n3786), .Y(n479) );
  OAI221XL U4587 ( .A0(n4019), .A1(n478), .B0(n1587), .B1(n4045), .C0(n482), 
        .Y(n2621) );
  AOI22X1 U4588 ( .A0(N262), .A1(n3790), .B0(N1001), .B1(n3786), .Y(n482) );
  OAI221XL U4589 ( .A0(n4020), .A1(n3783), .B0(n1588), .B1(n4045), .C0(n483), 
        .Y(n2622) );
  AOI22X1 U4590 ( .A0(N261), .A1(n3790), .B0(N1000), .B1(n3786), .Y(n483) );
  OAI221XL U4591 ( .A0(n4021), .A1(n478), .B0(n1589), .B1(n4045), .C0(n484), 
        .Y(n2623) );
  AOI22X1 U4592 ( .A0(N260), .A1(n3790), .B0(N999), .B1(n3786), .Y(n484) );
  OAI221XL U4593 ( .A0(n4022), .A1(n3783), .B0(n1590), .B1(n4045), .C0(n485), 
        .Y(n2624) );
  AOI22X1 U4594 ( .A0(N259), .A1(n3790), .B0(N998), .B1(n3786), .Y(n485) );
  OAI221XL U4595 ( .A0(n2686), .A1(n478), .B0(n1591), .B1(n4045), .C0(n486), 
        .Y(n2625) );
  AOI22X1 U4596 ( .A0(N258), .A1(n3790), .B0(N997), .B1(n3786), .Y(n486) );
  OAI221XL U4597 ( .A0(n2693), .A1(n3783), .B0(n1592), .B1(n4045), .C0(n487), 
        .Y(n2626) );
  AOI22X1 U4598 ( .A0(N257), .A1(n3789), .B0(N996), .B1(n3786), .Y(n487) );
  OAI221XL U4599 ( .A0(n2683), .A1(n478), .B0(n1593), .B1(n4045), .C0(n490), 
        .Y(n2627) );
  AOI22X1 U4600 ( .A0(N256), .A1(n3789), .B0(N995), .B1(n3785), .Y(n490) );
  OAI221XL U4601 ( .A0(n4023), .A1(n3783), .B0(n1594), .B1(n4045), .C0(n501), 
        .Y(n2628) );
  AOI22X1 U4602 ( .A0(N255), .A1(n3788), .B0(N994), .B1(n3784), .Y(n501) );
  OAI221XL U4603 ( .A0(n4024), .A1(n478), .B0(n1595), .B1(n4045), .C0(n512), 
        .Y(n2629) );
  AOI22X1 U4604 ( .A0(N254), .A1(n3788), .B0(N993), .B1(n3784), .Y(n512) );
  NOR4X1 U4605 ( .A(n570), .B(n571), .C(n572), .D(n573), .Y(n564) );
  NOR4X1 U4606 ( .A(n566), .B(n567), .C(n568), .D(n569), .Y(n565) );
  NAND4X1 U4607 ( .A(n49), .B(n48), .C(n47), .D(n46), .Y(n570) );
  NOR2BX1 U4608 ( .AN(n213), .B(instruction[24]), .Y(n164) );
  NAND4X1 U4609 ( .A(n1605), .B(n1606), .C(counter[1]), .D(counter[0]), .Y(
        n566) );
  AND2X2 U4610 ( .A(instruction[24]), .B(n213), .Y(n179) );
  OAI221XL U4611 ( .A0(n4030), .A1(n238), .B0(N244), .B1(n3792), .C0(n240), 
        .Y(n234) );
  AOI221XL U4612 ( .A0(n3998), .A1(n4040), .B0(n242), .B1(instruction[9]), 
        .C0(n243), .Y(n240) );
  OAI221XL U4613 ( .A0(n4031), .A1(n3773), .B0(N245), .B1(n3792), .C0(n262), 
        .Y(n260) );
  AOI221XL U4614 ( .A0(n3998), .A1(n4041), .B0(n242), .B1(instruction[8]), 
        .C0(n243), .Y(n262) );
  OAI221XL U4615 ( .A0(n4034), .A1(n238), .B0(N248), .B1(n3792), .C0(n286), 
        .Y(n284) );
  AOI221XL U4616 ( .A0(n3998), .A1(n4044), .B0(n242), .B1(instruction[5]), 
        .C0(n243), .Y(n286) );
  OAI221XL U4617 ( .A0(n4033), .A1(n3773), .B0(N247), .B1(n3792), .C0(n278), 
        .Y(n276) );
  AOI221XL U4618 ( .A0(n3998), .A1(n4043), .B0(n242), .B1(instruction[6]), 
        .C0(n243), .Y(n278) );
  OAI221XL U4619 ( .A0(n4032), .A1(n238), .B0(N246), .B1(n3792), .C0(n270), 
        .Y(n268) );
  AOI221XL U4620 ( .A0(n3998), .A1(n4042), .B0(n242), .B1(instruction[7]), 
        .C0(n243), .Y(n270) );
  NAND4X1 U4621 ( .A(n45), .B(n44), .C(n43), .D(n42), .Y(n569) );
  NAND4X1 U4622 ( .A(n61), .B(n60), .C(n59), .D(n58), .Y(n573) );
  NAND4X1 U4623 ( .A(n41), .B(n40), .C(n1599), .D(n1600), .Y(n568) );
  NAND4X1 U4624 ( .A(n57), .B(n56), .C(n55), .D(n54), .Y(n572) );
  NAND4X1 U4625 ( .A(n1601), .B(n1602), .C(n1603), .D(n1604), .Y(n567) );
  NAND4X1 U4626 ( .A(n53), .B(n52), .C(n51), .D(n50), .Y(n571) );
  AND2X2 U4627 ( .A(N60), .B(n3973), .Y(N126) );
  NOR3X1 U4628 ( .A(n4004), .B(instruction[26]), .C(n4002), .Y(n553) );
  AND2X2 U4629 ( .A(instruction[21]), .B(instruction[20]), .Y(n154) );
  AND2X2 U4630 ( .A(instruction[21]), .B(n4007), .Y(n158) );
  NOR3X1 U4631 ( .A(instruction[26]), .B(instruction[27]), .C(n4004), .Y(n560)
         );
  NAND4X1 U4632 ( .A(instruction[26]), .B(instruction[25]), .C(n554), .D(n4002), .Y(n245) );
  NAND4X1 U4633 ( .A(instruction[27]), .B(n554), .C(n4004), .D(n4003), .Y(n476) );
  AND4X1 U4634 ( .A(n540), .B(instruction[29]), .C(instruction[30]), .D(n4001), 
        .Y(n536) );
  NOR3X1 U4635 ( .A(instruction[29]), .B(instruction[31]), .C(n4001), .Y(n563)
         );
  AND4X1 U4636 ( .A(instruction[31]), .B(n553), .C(n552), .D(n3999), .Y(n3778)
         );
  CLKINVX1 U4637 ( .A(instruction[25]), .Y(n4004) );
  AND4X1 U4638 ( .A(instruction[31]), .B(n553), .C(n552), .D(n3999), .Y(n251)
         );
  AND4X1 U4639 ( .A(n551), .B(instruction[31]), .C(n552), .D(n3999), .Y(n3782)
         );
  AND4X1 U4640 ( .A(n551), .B(instruction[31]), .C(n552), .D(n3999), .Y(n249)
         );
  AND4X1 U4641 ( .A(n540), .B(instruction[28]), .C(n4000), .D(n3999), .Y(n518)
         );
  AND2X2 U4642 ( .A(n525), .B(instruction[31]), .Y(n540) );
  AND2X2 U4643 ( .A(n563), .B(instruction[30]), .Y(n561) );
  AND4X1 U4644 ( .A(instruction[27]), .B(instruction[26]), .C(n554), .D(n4004), 
        .Y(n3776) );
  AND4X1 U4645 ( .A(instruction[27]), .B(instruction[26]), .C(n554), .D(n4004), 
        .Y(n3775) );
  AND4X1 U4646 ( .A(instruction[27]), .B(instruction[26]), .C(n554), .D(n4004), 
        .Y(n254) );
  NOR2X1 U4647 ( .A(n4005), .B(instruction[22]), .Y(n190) );
  NOR2X1 U4648 ( .A(instruction[22]), .B(instruction[23]), .Y(n203) );
  NOR2X1 U4649 ( .A(n4006), .B(instruction[23]), .Y(n163) );
  AND4X1 U4650 ( .A(n540), .B(instruction[28]), .C(instruction[30]), .D(n4000), 
        .Y(n516) );
  AND2X2 U4651 ( .A(n539), .B(instruction[30]), .Y(n515) );
  CLKINVX1 U4652 ( .A(n545), .Y(n3995) );
  OAI211X1 U4653 ( .A0(instruction[31]), .A1(instruction[30]), .B0(n546), .C0(
        n525), .Y(n545) );
  OAI21XL U4654 ( .A0(instruction[28]), .A1(n3999), .B0(instruction[29]), .Y(
        n546) );
  AND3X2 U4655 ( .A(n553), .B(n543), .C(instruction[31]), .Y(n470) );
  CLKINVX1 U4656 ( .A(instruction[26]), .Y(n4003) );
  CLKINVX1 U4657 ( .A(instruction[27]), .Y(n4002) );
  CLKINVX1 U4658 ( .A(instruction[9]), .Y(n4040) );
  CLKINVX1 U4659 ( .A(instruction[8]), .Y(n4041) );
  CLKINVX1 U4660 ( .A(instruction[7]), .Y(n4042) );
  CLKINVX1 U4661 ( .A(instruction[6]), .Y(n4043) );
  CLKINVX1 U4662 ( .A(instruction[5]), .Y(n4044) );
  CLKINVX1 U4663 ( .A(instruction[22]), .Y(n4006) );
  CLKINVX1 U4664 ( .A(instruction[23]), .Y(n4005) );
  CLKINVX1 U4665 ( .A(instruction[20]), .Y(n4007) );
  CLKINVX1 U4666 ( .A(instruction[29]), .Y(n4000) );
  AND2X1 U4667 ( .A(\sub_1_root_add_0_root_add_137_ni_b0/carry[13] ), .B(n3978), .Y(\sub_1_root_add_0_root_add_137_ni_b0/carry[14] ) );
  XOR2X1 U4668 ( .A(n3978), .B(\sub_1_root_add_0_root_add_137_ni_b0/carry[13] ), .Y(N643) );
  AND2X1 U4669 ( .A(\sub_1_root_add_0_root_add_137_ni_b0/carry[12] ), .B(n3979), .Y(\sub_1_root_add_0_root_add_137_ni_b0/carry[13] ) );
  XOR2X1 U4670 ( .A(n3979), .B(\sub_1_root_add_0_root_add_137_ni_b0/carry[12] ), .Y(N644) );
  AND2X1 U4671 ( .A(\sub_1_root_add_0_root_add_137_ni_b0/carry[11] ), .B(n3981), .Y(\sub_1_root_add_0_root_add_137_ni_b0/carry[12] ) );
  XOR2X1 U4672 ( .A(n3981), .B(\sub_1_root_add_0_root_add_137_ni_b0/carry[11] ), .Y(N645) );
  AND2X1 U4673 ( .A(\sub_1_root_add_0_root_add_137_ni_b0/carry[10] ), .B(n3982), .Y(\sub_1_root_add_0_root_add_137_ni_b0/carry[11] ) );
  XOR2X1 U4674 ( .A(n3982), .B(\sub_1_root_add_0_root_add_137_ni_b0/carry[10] ), .Y(N646) );
  AND2X1 U4675 ( .A(\sub_1_root_add_0_root_add_137_ni_b0/carry[9] ), .B(n4040), 
        .Y(\sub_1_root_add_0_root_add_137_ni_b0/carry[10] ) );
  XOR2X1 U4676 ( .A(n4040), .B(\sub_1_root_add_0_root_add_137_ni_b0/carry[9] ), 
        .Y(N647) );
  AND2X1 U4677 ( .A(\sub_1_root_add_0_root_add_137_ni_b0/carry[8] ), .B(n4041), 
        .Y(\sub_1_root_add_0_root_add_137_ni_b0/carry[9] ) );
  XOR2X1 U4678 ( .A(n4041), .B(\sub_1_root_add_0_root_add_137_ni_b0/carry[8] ), 
        .Y(N648) );
  AND2X1 U4679 ( .A(\sub_1_root_add_0_root_add_137_ni_b0/carry[7] ), .B(n4042), 
        .Y(\sub_1_root_add_0_root_add_137_ni_b0/carry[8] ) );
  XOR2X1 U4680 ( .A(n4042), .B(\sub_1_root_add_0_root_add_137_ni_b0/carry[7] ), 
        .Y(N649) );
  AND2X1 U4681 ( .A(\sub_1_root_add_0_root_add_137_ni_b0/carry[6] ), .B(n4043), 
        .Y(\sub_1_root_add_0_root_add_137_ni_b0/carry[7] ) );
  AND2X1 U4682 ( .A(\sub_1_root_add_0_root_add_137_ni_b0/carry[5] ), .B(n4044), 
        .Y(\sub_1_root_add_0_root_add_137_ni_b0/carry[6] ) );
  XOR2X1 U4683 ( .A(n4044), .B(\sub_1_root_add_0_root_add_137_ni_b0/carry[5] ), 
        .Y(N651) );
  AND2X1 U4684 ( .A(\sub_1_root_add_0_root_add_137_ni_b0/carry[4] ), .B(n3977), 
        .Y(\sub_1_root_add_0_root_add_137_ni_b0/carry[5] ) );
  XOR2X1 U4685 ( .A(n3977), .B(\sub_1_root_add_0_root_add_137_ni_b0/carry[4] ), 
        .Y(N652) );
  AND2X1 U4686 ( .A(\sub_1_root_add_0_root_add_137_ni_b0/carry[3] ), .B(n3976), 
        .Y(\sub_1_root_add_0_root_add_137_ni_b0/carry[4] ) );
  XOR2X1 U4687 ( .A(n3976), .B(\sub_1_root_add_0_root_add_137_ni_b0/carry[3] ), 
        .Y(N653) );
  AND2X1 U4688 ( .A(\sub_1_root_add_0_root_add_137_ni_b0/carry[2] ), .B(n3975), 
        .Y(\sub_1_root_add_0_root_add_137_ni_b0/carry[3] ) );
  XOR2X1 U4689 ( .A(n3975), .B(\sub_1_root_add_0_root_add_137_ni_b0/carry[2] ), 
        .Y(N654) );
  AND2X1 U4690 ( .A(n3787), .B(n3974), .Y(
        \sub_1_root_add_0_root_add_137_ni_b0/carry[2] ) );
  XOR2X1 U4691 ( .A(n3974), .B(n3787), .Y(N655) );
  XNOR2X1 U4692 ( .A(\seIM[31] ), .B(
        \sub_1_root_add_0_root_add_137_ni_b0/carry[14] ), .Y(N642) );
  NOR4X1 U4693 ( .A(counter[27]), .B(counter[26]), .C(counter[25]), .D(
        counter[24]), .Y(n3986) );
  NOR4X1 U4694 ( .A(counter[30]), .B(counter[2]), .C(counter[29]), .D(
        counter[28]), .Y(n3985) );
  NOR4X1 U4695 ( .A(counter[5]), .B(counter[4]), .C(counter[3]), .D(
        counter[31]), .Y(n3984) );
  NOR4X1 U4696 ( .A(counter[9]), .B(counter[8]), .C(counter[7]), .D(counter[6]), .Y(n3983) );
  NAND4X1 U4697 ( .A(n3986), .B(n3985), .C(n3984), .D(n3983), .Y(n3992) );
  AOI211X1 U4698 ( .A0(counter[1]), .A1(counter[0]), .B0(counter[11]), .C0(
        counter[10]), .Y(n3990) );
  NOR4X1 U4699 ( .A(counter[15]), .B(counter[14]), .C(counter[13]), .D(
        counter[12]), .Y(n3989) );
  NOR4X1 U4700 ( .A(counter[19]), .B(counter[18]), .C(counter[17]), .D(
        counter[16]), .Y(n3988) );
  NOR4X1 U4701 ( .A(counter[23]), .B(counter[22]), .C(counter[21]), .D(
        counter[20]), .Y(n3987) );
  NAND4X1 U4702 ( .A(n3990), .B(n3989), .C(n3988), .D(n3987), .Y(n3991) );
endmodule

