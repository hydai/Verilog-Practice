`timescale 1ns / 1ps

module display_ctrl(pattern, reset, clk, startStop, Pause);
	parameter INIT = 2'd0;
	parameter RUN = 2'd1;
	parameter PAUSE = 2'd2;
	input clk;
	input reset;
	input startStop, Pause;
	output [255:0] pattern;
	integer ct;
	wire startStop_op, Pause_op;
	reg [255:0] pattern;
	reg [3:0] state;
	reg [255:0] graph [12:0];
	// Get LGS
	always @(*) begin
		pattern = graph[ct];
	end
	
	one_pulse op1(startStop_op, !startStop, clk, reset);
	one_pulse op2(Pause_op, !Pause, clk, reset);
	
	// Store state
	always @(posedge clk or negedge reset) begin
		if (!reset) begin
			state <= INIT;
			ct <= 0;
		end else if (Pause_op) begin
			if (state == INIT) begin
				state <= INIT;
				ct <= 0;
			end else begin
				state <= PAUSE;
				ct <= ct;
			end
		end else if (startStop_op) begin
			if (state == INIT) begin
				state <= RUN;
				ct <= ct;
			end else if (state == RUN) begin
				state <= INIT;
				ct <= 0;
			end else begin
				state <= RUN;
				ct <= ct;
			end
		end else if (state == RUN) begin
			state <= state;
			if (ct + 1'b1 > 12) begin
				ct <= 1'b1;
			end else begin
				ct <= ct + 1'b1;
			end
		end else begin
			state <= state;
			ct <= ct;
		end
	end

	always @(*) begin
		 graph[0] = 256'b0000000000000000000000000000000000000000000000000000111111110000000010000001000000000100001000000000001001000000000000011000000000000001100000000000001001000000000001000010000000001000000100000000111111110000000000000000000000000000000000000000000000000000;
		 graph[1] = 256'b0000000000000000000000000000000000000000000000000000111111110000000011111111000000000111111000000000001111000000000000011000000000000001100000000000001001000000000001000010000000001000000100000000111111110000000000000000000000000000000000000000000000000000;
		 graph[2] = 256'b0000000000000000000000000000000000000000000000000000111111110000000010111101000000000111111000000000001111000000000000011000000000000001100000000000001001000000000001000010000000001001100100000000111111110000000000000000000000000000000000000000000000000000;
		 graph[3] = 256'b0000000000000000000000000000000000000000000000000000111111110000000010011001000000000111111000000000001111000000000000011000000000000001100000000000001001000000000001000010000000001011110100000000111111110000000000000000000000000000000000000000000000000000;
		 graph[4] = 256'b0000000000000000000000000000000000000000000000000000111111110000000010000001000000000111111000000000001111000000000000011000000000000001100000000000001001000000000001000010000000001111111100000000111111110000000000000000000000000000000000000000000000000000;
		 graph[5] = 256'b0000000000000000000000000000000000000000000000000000111111110000000010000001000000000101101000000000001111000000000000011000000000000001100000000000001001000000000001011010000000001111111100000000111111110000000000000000000000000000000000000000000000000000;
		 graph[6] = 256'b0000000000000000000000000000000000000000000000000000111111110000000010000001000000000100001000000000001111000000000000011000000000000001100000000000001001000000000001111110000000001111111100000000111111110000000000000000000000000000000000000000000000000000;
		 graph[7] = 256'b0000000000000000000000000000000000000000000000000000111111110000000010000001000000000100001000000000001001000000000000011000000000000001100000000000001111000000000001111110000000001111111100000000111111110000000000000000000000000000000000000000000000000000;
		 graph[8] = 256'b0000000000000000000000000000000000000111000000000000011111110000000001000111100000000010001110000000001101110000000000011100000000000011100000000000011111000000000111111110000000011111111000000000011111100000000000000110000000000000000000000000000000000000;
		 graph[9] = 256'b0000000000000000000000000000000000000011100000000000001011100000000000010011000000000001000111000000000100011100000000011111000000001111100000000011111110000000001111111000000000001111110000000000001111100000000000001110000000000000000000000000000000000000;
		 graph[10] = 256'b0000000000000000000000000000000000000000000000000000000000000000000110000001100000010100001010000001001001001000000100011000100000010001100010000001001001001000000101000010100000011000000110000000000000000000000000000000000000000000000000000000000000000000;
		 graph[11] = 256'b0000000000000000000000000000000000000000000000000000110000000000000011100000000000001110000011000001111101111100000111111100110000011111100010000011111010001000001100000101100000000000010100000000000000110000000000000001000000000000000000000000000000000000;
		 graph[12] = 256'b000000000000000000000000000000000000001100000000000001110000000000011111000000000011111100000000011111110000000001111111011010000111001101101000000000010001100000000001001100000000000101100000000000011100000000000001100000000000000000000000000000000000000;
	end

endmodule

/*
	assign LGS[15*16+:16] = 16'b0000_0011_1000_0000;
	assign LGS[14*16+:16] = 16'b0000_0011_1000_0000;
	assign LGS[13*16+:16] = 16'b0000_0011_1000_0000;
	assign LGS[12*16+:16] = 16'b0000_0010_1000_0000;
	assign LGS[11*16+:16] = 16'b0000_0111_1100_0000;
	assign LGS[10*16+:16] = 16'b0000_1111_1110_0000;
	assign LGS[ 9*16+:16] = 16'b0001_1111_1111_0000;
	assign LGS[ 8*16+:16] = 16'b0001_1011_1011_0000;
	assign LGS[ 7*16+:16] = 16'b0001_1011_1011_0000;
	assign LGS[ 6*16+:16] = 16'b0001_1011_1011_0000;
	assign LGS[ 5*16+:16] = 16'b0001_0111_1101_0000;
	assign LGS[ 4*16+:16] = 16'b0000_0110_1100_0000;
	assign LGS[ 3*16+:16] = 16'b0000_0110_1100_0000;
	assign LGS[ 2*16+:16] = 16'b0000_0110_1100_0000;
	assign LGS[ 1*16+:16] = 16'b0000_1110_1110_0000;
	assign LGS[ 0*16+:16] = 16'b0001_1110_1111_0000;
	*/