
module datapath_DW01_inc_0 ( A, SUM );
  input [16:0] A;
  output [16:0] SUM;

  wire   [16:2] carry;

  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXL U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(SUM[16]), .S(SUM[15]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module datapath_DW_rightsh_1 ( A, DATA_TC, SH, B );
  input [15:0] A;
  input [31:0] SH;
  output [15:0] B;
  input DATA_TC;
  wire   n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235;

  OR2XL U128 ( .A(n226), .B(SH[2]), .Y(n195) );
  MX2XL U129 ( .A(n202), .B(n223), .S0(SH[2]), .Y(n190) );
  MXI2XL U130 ( .A(n198), .B(n227), .S0(SH[2]), .Y(n217) );
  MXI2XL U131 ( .A(n194), .B(n226), .S0(SH[2]), .Y(n210) );
  OR2XL U132 ( .A(n223), .B(SH[2]), .Y(n203) );
  OR2XL U133 ( .A(n230), .B(SH[2]), .Y(n207) );
  MX3X1 U134 ( .A(n235), .B(n187), .C(n191), .S0(SH[2]), .S1(n182), .Y(n234)
         );
  MX3X1 U135 ( .A(n211), .B(n212), .C(n179), .S0(n189), .S1(SH[2]), .Y(n209)
         );
  CLKMX2X2 U136 ( .A(A[7]), .B(A[8]), .S0(n183), .Y(n214) );
  CLKMX2X2 U137 ( .A(A[10]), .B(A[11]), .S0(n183), .Y(n233) );
  NOR2X1 U138 ( .A(n215), .B(n181), .Y(B[2]) );
  CLKINVX1 U139 ( .A(SH[1]), .Y(n189) );
  CLKINVX1 U140 ( .A(n234), .Y(n185) );
  NOR2XL U141 ( .A(n180), .B(n185), .Y(B[0]) );
  MXI2X1 U142 ( .A(n209), .B(n210), .S0(n182), .Y(n208) );
  NOR2X1 U143 ( .A(n196), .B(n180), .Y(B[6]) );
  INVXL U144 ( .A(n225), .Y(n186) );
  CLKMX2X2 U145 ( .A(n213), .B(n214), .S0(n189), .Y(n179) );
  MXI2XL U146 ( .A(n213), .B(n214), .S0(n189), .Y(n193) );
  NOR3XL U147 ( .A(n190), .B(n180), .C(n182), .Y(B[9]) );
  NOR3XL U148 ( .A(n203), .B(n180), .C(n182), .Y(B[13]) );
  NOR3XL U149 ( .A(n199), .B(n180), .C(n182), .Y(B[14]) );
  NOR3XL U150 ( .A(n195), .B(n180), .C(n182), .Y(B[15]) );
  NOR3XL U151 ( .A(n207), .B(n180), .C(n182), .Y(B[12]) );
  OR2XL U152 ( .A(n227), .B(SH[2]), .Y(n199) );
  CLKINVX1 U153 ( .A(n197), .Y(n188) );
  CLKINVX1 U154 ( .A(n205), .Y(n187) );
  NOR3BXL U155 ( .AN(n191), .B(n180), .C(n182), .Y(B[8]) );
  CLKBUFX3 U156 ( .A(SH[4]), .Y(n180) );
  NOR3BXL U157 ( .AN(n217), .B(n180), .C(n182), .Y(B[10]) );
  NOR3BXL U158 ( .AN(n210), .B(n180), .C(n182), .Y(B[11]) );
  CLKBUFX3 U159 ( .A(SH[4]), .Y(n181) );
  NOR2X1 U160 ( .A(n200), .B(n180), .Y(B[5]) );
  NOR2X1 U161 ( .A(n204), .B(n181), .Y(B[4]) );
  NOR2X1 U162 ( .A(n208), .B(n181), .Y(B[3]) );
  NOR2X1 U163 ( .A(n192), .B(n180), .Y(B[7]) );
  NOR2X1 U164 ( .A(n222), .B(n180), .Y(B[1]) );
  CLKBUFX3 U165 ( .A(SH[0]), .Y(n183) );
  CLKBUFX3 U166 ( .A(SH[0]), .Y(n184) );
  CLKBUFX3 U167 ( .A(SH[3]), .Y(n182) );
  MX3XL U168 ( .A(n193), .B(n194), .C(n195), .S0(SH[2]), .S1(n182), .Y(n192)
         );
  MX3XL U169 ( .A(n197), .B(n198), .C(n199), .S0(SH[2]), .S1(n182), .Y(n196)
         );
  MX3XL U170 ( .A(n201), .B(n202), .C(n203), .S0(SH[2]), .S1(n182), .Y(n200)
         );
  MX3XL U171 ( .A(n205), .B(n206), .C(n207), .S0(SH[2]), .S1(n182), .Y(n204)
         );
  MXI2X1 U172 ( .A(n216), .B(n217), .S0(n182), .Y(n215) );
  MX3XL U173 ( .A(n218), .B(n219), .C(n188), .S0(n189), .S1(SH[2]), .Y(n216)
         );
  MXI2X1 U174 ( .A(n220), .B(n221), .S0(n189), .Y(n197) );
  MX3XL U175 ( .A(n186), .B(n201), .C(n190), .S0(SH[2]), .S1(n182), .Y(n222)
         );
  MXI2X1 U176 ( .A(n224), .B(n213), .S0(n189), .Y(n202) );
  CLKMX2X2 U177 ( .A(A[9]), .B(A[10]), .S0(n183), .Y(n213) );
  MXI2X1 U178 ( .A(n214), .B(n211), .S0(n189), .Y(n201) );
  CLKMX2X2 U179 ( .A(A[5]), .B(A[6]), .S0(n183), .Y(n211) );
  MX3XL U180 ( .A(A[1]), .B(A[2]), .C(n212), .S0(n184), .S1(SH[1]), .Y(n225)
         );
  CLKMX2X2 U181 ( .A(A[3]), .B(A[4]), .S0(n183), .Y(n212) );
  MXI2X1 U182 ( .A(n228), .B(n229), .S0(n189), .Y(n223) );
  NAND2X1 U183 ( .A(n228), .B(n189), .Y(n226) );
  NOR2BX1 U184 ( .AN(A[15]), .B(n184), .Y(n228) );
  MXI2X1 U185 ( .A(n229), .B(n224), .S0(n189), .Y(n194) );
  CLKMX2X2 U186 ( .A(A[11]), .B(A[12]), .S0(n183), .Y(n224) );
  CLKMX2X2 U187 ( .A(A[13]), .B(A[14]), .S0(n183), .Y(n229) );
  NAND2X1 U188 ( .A(n231), .B(n189), .Y(n227) );
  MXI2X1 U189 ( .A(n232), .B(n233), .S0(n189), .Y(n198) );
  MXI2X1 U190 ( .A(n206), .B(n230), .S0(SH[2]), .Y(n191) );
  MXI2X1 U191 ( .A(n231), .B(n232), .S0(n189), .Y(n230) );
  CLKMX2X2 U192 ( .A(A[12]), .B(A[13]), .S0(n183), .Y(n232) );
  CLKMX2X2 U193 ( .A(A[14]), .B(A[15]), .S0(n183), .Y(n231) );
  MXI2X1 U194 ( .A(n233), .B(n220), .S0(n189), .Y(n206) );
  CLKMX2X2 U195 ( .A(A[8]), .B(A[9]), .S0(n183), .Y(n220) );
  MXI2X1 U196 ( .A(n221), .B(n218), .S0(n189), .Y(n205) );
  CLKMX2X2 U197 ( .A(A[4]), .B(A[5]), .S0(n183), .Y(n218) );
  CLKMX2X2 U198 ( .A(A[6]), .B(A[7]), .S0(n183), .Y(n221) );
  MX3XL U199 ( .A(A[0]), .B(A[1]), .C(n219), .S0(n184), .S1(SH[1]), .Y(n235)
         );
  CLKMX2X2 U200 ( .A(A[2]), .B(A[3]), .S0(n183), .Y(n219) );
endmodule


module datapath_DW_leftsh_0 ( A, SH, B );
  input [15:0] A;
  input [31:0] SH;
  output [15:0] B;
  wire   n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233;

  INVX3 U127 ( .A(SH[2]), .Y(n182) );
  INVX1 U128 ( .A(SH[1]), .Y(n187) );
  MXI2X1 U129 ( .A(n226), .B(n227), .S0(n187), .Y(n193) );
  MXI2X1 U130 ( .A(n219), .B(n217), .S0(n187), .Y(n205) );
  MXI2X1 U131 ( .A(n218), .B(n221), .S0(n187), .Y(n206) );
  NOR3X1 U132 ( .A(n195), .B(n177), .C(n179), .Y(B[0]) );
  NAND2BX1 U133 ( .AN(n202), .B(n182), .Y(n191) );
  MX2XL U134 ( .A(n211), .B(n212), .S0(SH[2]), .Y(n197) );
  MXI2XL U135 ( .A(n227), .B(n229), .S0(n187), .Y(n211) );
  MXI2XL U136 ( .A(n222), .B(n220), .S0(n187), .Y(n208) );
  MXI2XL U137 ( .A(n230), .B(n228), .S0(n187), .Y(n210) );
  MXI2XL U138 ( .A(n205), .B(n206), .S0(n182), .Y(n196) );
  NAND2XL U139 ( .A(n219), .B(n187), .Y(n202) );
  INVXL U140 ( .A(n190), .Y(n186) );
  INVXL U141 ( .A(n194), .Y(n185) );
  AND2XL U142 ( .A(A[0]), .B(n180), .Y(n233) );
  MX2XL U143 ( .A(A[11]), .B(A[10]), .S0(SH[0]), .Y(n220) );
  CLKINVX1 U144 ( .A(n208), .Y(n184) );
  NOR3X1 U145 ( .A(n201), .B(n177), .C(n179), .Y(B[2]) );
  NOR3X1 U146 ( .A(n191), .B(n177), .C(n179), .Y(B[1]) );
  NOR3X1 U147 ( .A(n200), .B(n177), .C(n179), .Y(B[3]) );
  NOR3X1 U148 ( .A(n197), .B(n177), .C(n179), .Y(B[6]) );
  NOR3BXL U149 ( .AN(n199), .B(n177), .C(n179), .Y(B[4]) );
  NOR3BXL U150 ( .AN(n198), .B(n177), .C(n179), .Y(B[5]) );
  NOR3BXL U151 ( .AN(n196), .B(n177), .C(n179), .Y(B[7]) );
  CLKBUFX3 U152 ( .A(SH[4]), .Y(n177) );
  CLKBUFX3 U153 ( .A(SH[4]), .Y(n178) );
  NOR2X1 U154 ( .A(n223), .B(n177), .Y(B[12]) );
  NOR2X1 U155 ( .A(n209), .B(n177), .Y(B[14]) );
  CLKINVX1 U156 ( .A(n213), .Y(n183) );
  NOR2X1 U157 ( .A(n192), .B(n178), .Y(B[8]) );
  NOR2X1 U158 ( .A(n188), .B(n177), .Y(B[9]) );
  NOR2X1 U159 ( .A(n232), .B(n178), .Y(B[10]) );
  NOR2X1 U160 ( .A(n215), .B(n177), .Y(B[13]) );
  CLKBUFX3 U161 ( .A(SH[3]), .Y(n179) );
  NOR2X1 U162 ( .A(n177), .B(n181), .Y(B[15]) );
  CLKINVX1 U163 ( .A(n203), .Y(n181) );
  CLKINVX1 U164 ( .A(SH[0]), .Y(n180) );
  NOR2X1 U165 ( .A(n231), .B(n178), .Y(B[11]) );
  MX3XL U166 ( .A(n189), .B(n190), .C(n191), .S0(n182), .S1(n179), .Y(n188) );
  MX3XL U167 ( .A(n193), .B(n194), .C(n195), .S0(n182), .S1(n179), .Y(n192) );
  MX3XL U168 ( .A(n184), .B(n204), .C(n196), .S0(n182), .S1(n179), .Y(n203) );
  MX3XL U169 ( .A(A[14]), .B(A[15]), .C(n207), .S0(n180), .S1(SH[1]), .Y(n204)
         );
  MX3XL U170 ( .A(n210), .B(n183), .C(n197), .S0(n182), .S1(n179), .Y(n209) );
  MX3XL U171 ( .A(A[13]), .B(A[14]), .C(n214), .S0(n180), .S1(SH[1]), .Y(n213)
         );
  MXI2X1 U172 ( .A(n216), .B(n198), .S0(n179), .Y(n215) );
  MXI2X1 U173 ( .A(n202), .B(n189), .S0(n182), .Y(n198) );
  MXI2X1 U174 ( .A(n217), .B(n218), .S0(n187), .Y(n189) );
  MX3XL U175 ( .A(n220), .B(n207), .C(n186), .S0(n187), .S1(SH[2]), .Y(n216)
         );
  MXI2X1 U176 ( .A(n221), .B(n222), .S0(n187), .Y(n190) );
  CLKMX2X2 U177 ( .A(A[13]), .B(A[12]), .S0(SH[0]), .Y(n207) );
  MXI2X1 U178 ( .A(n224), .B(n199), .S0(n179), .Y(n223) );
  MXI2X1 U179 ( .A(n225), .B(n193), .S0(n182), .Y(n199) );
  MX3XL U180 ( .A(n228), .B(n214), .C(n185), .S0(n187), .S1(SH[2]), .Y(n224)
         );
  MXI2X1 U181 ( .A(n229), .B(n230), .S0(n187), .Y(n194) );
  CLKMX2X2 U182 ( .A(A[12]), .B(A[11]), .S0(SH[0]), .Y(n214) );
  MX3XL U183 ( .A(n206), .B(n208), .C(n200), .S0(n182), .S1(n179), .Y(n231) );
  NAND2BX1 U184 ( .AN(n205), .B(n182), .Y(n200) );
  CLKMX2X2 U185 ( .A(A[3]), .B(A[2]), .S0(SH[0]), .Y(n217) );
  CLKMX2X2 U186 ( .A(A[1]), .B(A[0]), .S0(SH[0]), .Y(n219) );
  CLKMX2X2 U187 ( .A(A[9]), .B(A[8]), .S0(SH[0]), .Y(n222) );
  CLKMX2X2 U188 ( .A(A[7]), .B(A[6]), .S0(SH[0]), .Y(n221) );
  CLKMX2X2 U189 ( .A(A[5]), .B(A[4]), .S0(SH[0]), .Y(n218) );
  MX3XL U190 ( .A(n211), .B(n210), .C(n201), .S0(n182), .S1(n179), .Y(n232) );
  NAND2BX1 U191 ( .AN(n212), .B(n182), .Y(n201) );
  MXI2X1 U192 ( .A(n233), .B(n226), .S0(n187), .Y(n212) );
  CLKMX2X2 U193 ( .A(A[2]), .B(A[1]), .S0(SH[0]), .Y(n226) );
  CLKMX2X2 U194 ( .A(A[10]), .B(A[9]), .S0(SH[0]), .Y(n228) );
  CLKMX2X2 U195 ( .A(A[8]), .B(A[7]), .S0(SH[0]), .Y(n230) );
  CLKMX2X2 U196 ( .A(A[6]), .B(A[5]), .S0(SH[0]), .Y(n229) );
  CLKMX2X2 U197 ( .A(A[4]), .B(A[3]), .S0(SH[0]), .Y(n227) );
  NAND2BX1 U198 ( .AN(n225), .B(n182), .Y(n195) );
  NAND2X1 U199 ( .A(n233), .B(n187), .Y(n225) );
endmodule


module datapath_DW01_add_5 ( A, B, CI, SUM, CO );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n21, n23, n24, n25, n26, n27, n29, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n74, n76, n77, n78, n79, n80,
         n81, n84, n85, n86, n87, n88, n89, n94, n96, n99, n100, n163, n164,
         n165, n166, n167, n168, n169, n170, n171;

  XOR2X1 U16 ( .A(n27), .B(n3), .Y(SUM[13]) );
  XOR2X1 U30 ( .A(n35), .B(n5), .Y(SUM[11]) );
  XOR2X1 U44 ( .A(n43), .B(n7), .Y(SUM[9]) );
  XOR2X1 U61 ( .A(n54), .B(n9), .Y(SUM[7]) );
  XOR2X1 U67 ( .A(n59), .B(n10), .Y(SUM[6]) );
  XOR2X1 U102 ( .A(n84), .B(n14), .Y(SUM[2]) );
  XOR2X1 U112 ( .A(n15), .B(n88), .Y(SUM[1]) );
  OR2XL U125 ( .A(B[3]), .B(A[3]), .Y(n170) );
  INVX1 U126 ( .A(n35), .Y(n163) );
  OAI21XL U127 ( .A0(n72), .A1(n68), .B0(n69), .Y(n67) );
  NAND2X1 U128 ( .A(n163), .B(n164), .Y(n165) );
  NAND2X1 U129 ( .A(n165), .B(n34), .Y(n32) );
  NAND2X1 U130 ( .A(n166), .B(n167), .Y(n168) );
  NAND2X1 U131 ( .A(n168), .B(n87), .Y(n85) );
  CLKINVX1 U132 ( .A(n86), .Y(n166) );
  CLKINVX1 U133 ( .A(n88), .Y(n167) );
  NAND2X1 U134 ( .A(B[11]), .B(A[11]), .Y(n34) );
  NAND2X1 U135 ( .A(B[1]), .B(A[1]), .Y(n87) );
  NOR2X1 U136 ( .A(B[11]), .B(A[11]), .Y(n33) );
  CLKINVX1 U137 ( .A(n33), .Y(n164) );
  AOI21X1 U138 ( .A0(n32), .A1(n169), .B0(n29), .Y(n27) );
  INVXL U139 ( .A(n85), .Y(n84) );
  AOI21X1 U140 ( .A0(n85), .A1(n66), .B0(n67), .Y(n65) );
  NOR2X1 U141 ( .A(B[4]), .B(A[4]), .Y(n68) );
  INVXL U142 ( .A(n44), .Y(n43) );
  NOR2X1 U143 ( .A(n62), .B(n57), .Y(n55) );
  OAI21XL U144 ( .A0(n19), .A1(n17), .B0(n18), .Y(SUM[16]) );
  NAND2BXL U145 ( .AN(n86), .B(n87), .Y(n15) );
  NOR2X1 U146 ( .A(B[2]), .B(A[2]), .Y(n78) );
  NOR2XL U147 ( .A(B[1]), .B(A[1]), .Y(n86) );
  AOI21XL U148 ( .A0(n64), .A1(n55), .B0(n56), .Y(n54) );
  NAND2XL U149 ( .A(n170), .B(n76), .Y(n13) );
  NAND2BX1 U150 ( .AN(n25), .B(n26), .Y(n3) );
  NAND2BX1 U151 ( .AN(n33), .B(n34), .Y(n5) );
  NAND2BX1 U152 ( .AN(n41), .B(n42), .Y(n7) );
  INVXL U153 ( .A(n17), .Y(n89) );
  NAND2XL U154 ( .A(n80), .B(n79), .Y(n14) );
  NAND2BXL U155 ( .AN(n52), .B(n53), .Y(n9) );
  XNOR2XL U156 ( .A(n24), .B(n2), .Y(SUM[14]) );
  XNOR2XL U157 ( .A(n32), .B(n4), .Y(SUM[12]) );
  XNOR2XL U158 ( .A(n40), .B(n6), .Y(SUM[10]) );
  NAND2XL U159 ( .A(n99), .B(n63), .Y(n11) );
  INVXL U160 ( .A(n49), .Y(n96) );
  AOI21XL U161 ( .A0(n24), .A1(n171), .B0(n21), .Y(n19) );
  AOI21XL U162 ( .A0(n44), .A1(n36), .B0(n37), .Y(n35) );
  NAND2BXL U163 ( .AN(n57), .B(n58), .Y(n10) );
  NAND2XL U164 ( .A(n170), .B(n80), .Y(n71) );
  INVXL U165 ( .A(n63), .Y(n61) );
  NOR2XL U166 ( .A(B[0]), .B(A[0]), .Y(n88) );
  NOR2XL U167 ( .A(B[5]), .B(A[5]), .Y(n62) );
  NAND2XL U168 ( .A(B[3]), .B(A[3]), .Y(n76) );
  NAND2XL U169 ( .A(B[8]), .B(A[8]), .Y(n50) );
  NAND2XL U170 ( .A(B[4]), .B(A[4]), .Y(n69) );
  NAND2XL U171 ( .A(B[6]), .B(A[6]), .Y(n58) );
  XNOR2XL U172 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  CLKINVX1 U173 ( .A(n65), .Y(n64) );
  AOI21X1 U174 ( .A0(n64), .A1(n99), .B0(n61), .Y(n59) );
  OAI21XL U175 ( .A0(n65), .A1(n45), .B0(n46), .Y(n44) );
  NAND2X1 U176 ( .A(n55), .B(n47), .Y(n45) );
  AOI21X1 U177 ( .A0(n56), .A1(n47), .B0(n48), .Y(n46) );
  NOR2X1 U178 ( .A(n52), .B(n49), .Y(n47) );
  NOR2X1 U179 ( .A(n71), .B(n68), .Y(n66) );
  XNOR2X1 U180 ( .A(n51), .B(n8), .Y(SUM[8]) );
  NAND2X1 U181 ( .A(n96), .B(n50), .Y(n8) );
  OAI21XL U182 ( .A0(n54), .A1(n52), .B0(n53), .Y(n51) );
  NAND2X1 U183 ( .A(n94), .B(n39), .Y(n6) );
  OAI21XL U184 ( .A0(n43), .A1(n41), .B0(n42), .Y(n40) );
  CLKINVX1 U185 ( .A(n38), .Y(n94) );
  NAND2X1 U186 ( .A(n169), .B(n31), .Y(n4) );
  XNOR2X1 U187 ( .A(n77), .B(n13), .Y(SUM[3]) );
  OAI21XL U188 ( .A0(n84), .A1(n78), .B0(n79), .Y(n77) );
  XNOR2X1 U189 ( .A(n70), .B(n12), .Y(SUM[4]) );
  NAND2X1 U190 ( .A(n100), .B(n69), .Y(n12) );
  OAI21XL U191 ( .A0(n84), .A1(n71), .B0(n72), .Y(n70) );
  CLKINVX1 U192 ( .A(n68), .Y(n100) );
  XNOR2X1 U193 ( .A(n64), .B(n11), .Y(SUM[5]) );
  NAND2X1 U194 ( .A(n171), .B(n23), .Y(n2) );
  XOR2X1 U195 ( .A(n19), .B(n1), .Y(SUM[15]) );
  NAND2X1 U196 ( .A(n89), .B(n18), .Y(n1) );
  OAI21XL U197 ( .A0(n57), .A1(n63), .B0(n58), .Y(n56) );
  AOI21X1 U198 ( .A0(n170), .A1(n81), .B0(n74), .Y(n72) );
  CLKINVX1 U199 ( .A(n79), .Y(n81) );
  CLKINVX1 U200 ( .A(n76), .Y(n74) );
  OAI21XL U201 ( .A0(n27), .A1(n25), .B0(n26), .Y(n24) );
  CLKINVX1 U202 ( .A(n23), .Y(n21) );
  NOR2X1 U203 ( .A(n41), .B(n38), .Y(n36) );
  OAI21XL U204 ( .A0(n38), .A1(n42), .B0(n39), .Y(n37) );
  CLKINVX1 U205 ( .A(n31), .Y(n29) );
  OAI21XL U206 ( .A0(n49), .A1(n53), .B0(n50), .Y(n48) );
  CLKINVX1 U207 ( .A(n78), .Y(n80) );
  CLKINVX1 U208 ( .A(n62), .Y(n99) );
  NOR2X1 U209 ( .A(B[7]), .B(A[7]), .Y(n52) );
  NOR2X1 U210 ( .A(B[6]), .B(A[6]), .Y(n57) );
  NOR2X1 U211 ( .A(B[9]), .B(A[9]), .Y(n41) );
  NOR2X1 U212 ( .A(B[10]), .B(A[10]), .Y(n38) );
  NOR2X1 U213 ( .A(B[8]), .B(A[8]), .Y(n49) );
  NAND2X1 U214 ( .A(B[5]), .B(A[5]), .Y(n63) );
  NAND2X1 U215 ( .A(B[2]), .B(A[2]), .Y(n79) );
  NAND2X1 U216 ( .A(B[7]), .B(A[7]), .Y(n53) );
  NAND2X1 U217 ( .A(B[12]), .B(A[12]), .Y(n31) );
  NAND2X1 U218 ( .A(B[9]), .B(A[9]), .Y(n42) );
  OR2X1 U219 ( .A(B[12]), .B(A[12]), .Y(n169) );
  NAND2X1 U220 ( .A(B[10]), .B(A[10]), .Y(n39) );
  NOR2X1 U221 ( .A(B[13]), .B(A[13]), .Y(n25) );
  NOR2X1 U222 ( .A(B[15]), .B(A[15]), .Y(n17) );
  NAND2X1 U223 ( .A(B[14]), .B(A[14]), .Y(n23) );
  OR2X1 U224 ( .A(B[14]), .B(A[14]), .Y(n171) );
  NAND2X1 U225 ( .A(B[13]), .B(A[13]), .Y(n26) );
  NAND2X1 U226 ( .A(B[15]), .B(A[15]), .Y(n18) );
endmodule


module datapath_DW01_add_6 ( A, B, CI, SUM, CO );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n18, n19, n20, n22, n24, n25, n26, n27, n28, n30, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n75, n77, n78, n79, n80,
         n81, n82, n85, n86, n87, n88, n89, n90, n96, n97, n98, n102, n165,
         n166, n167, n168, n169, n170, n171;

  XOR2X1 U2 ( .A(n166), .B(n1), .Y(SUM[15]) );
  XOR2X1 U16 ( .A(n28), .B(n3), .Y(SUM[13]) );
  XOR2X1 U30 ( .A(n36), .B(n5), .Y(SUM[11]) );
  XOR2X1 U44 ( .A(n44), .B(n7), .Y(SUM[9]) );
  XOR2X1 U61 ( .A(n55), .B(n9), .Y(SUM[7]) );
  XOR2X1 U67 ( .A(n60), .B(n10), .Y(SUM[6]) );
  XOR2X1 U102 ( .A(n85), .B(n14), .Y(SUM[2]) );
  XOR2X1 U112 ( .A(n15), .B(n90), .Y(SUM[1]) );
  AOI21X1 U127 ( .A0(n25), .A1(n170), .B0(n22), .Y(n166) );
  OAI21X1 U128 ( .A0(n28), .A1(n26), .B0(n27), .Y(n25) );
  OAI21XL U129 ( .A0(n20), .A1(n18), .B0(n19), .Y(SUM[16]) );
  AND2X2 U130 ( .A(n56), .B(n48), .Y(n165) );
  OAI21XL U131 ( .A0(n87), .A1(n90), .B0(n88), .Y(n86) );
  NAND2XL U132 ( .A(B[0]), .B(A[0]), .Y(n90) );
  XNOR2XL U133 ( .A(n25), .B(n2), .Y(SUM[14]) );
  CLKINVX1 U134 ( .A(n66), .Y(n167) );
  AOI21X1 U135 ( .A0(n57), .A1(n48), .B0(n49), .Y(n47) );
  NAND2X1 U136 ( .A(n167), .B(n165), .Y(n168) );
  NAND2X1 U137 ( .A(n168), .B(n47), .Y(n45) );
  NAND2X1 U138 ( .A(B[5]), .B(A[5]), .Y(n64) );
  OR2X1 U139 ( .A(B[3]), .B(A[3]), .Y(n169) );
  OAI21XL U140 ( .A0(n73), .A1(n69), .B0(n70), .Y(n68) );
  NAND2BXL U141 ( .AN(n87), .B(n88), .Y(n15) );
  INVXL U142 ( .A(n39), .Y(n96) );
  NAND2BXL U143 ( .AN(n58), .B(n59), .Y(n10) );
  NOR2X1 U144 ( .A(B[8]), .B(A[8]), .Y(n50) );
  NOR2X1 U145 ( .A(B[7]), .B(A[7]), .Y(n53) );
  NOR2X1 U146 ( .A(B[6]), .B(A[6]), .Y(n58) );
  NAND2X1 U147 ( .A(B[7]), .B(A[7]), .Y(n54) );
  INVXL U148 ( .A(n45), .Y(n44) );
  AOI21XL U149 ( .A0(n65), .A1(n56), .B0(n57), .Y(n55) );
  NAND2BX1 U150 ( .AN(n18), .B(n19), .Y(n1) );
  NAND2BX1 U151 ( .AN(n26), .B(n27), .Y(n3) );
  NAND2XL U152 ( .A(n81), .B(n80), .Y(n14) );
  NAND2BX1 U153 ( .AN(n34), .B(n35), .Y(n5) );
  NAND2BX1 U154 ( .AN(n53), .B(n54), .Y(n9) );
  XNOR2XL U155 ( .A(n33), .B(n4), .Y(SUM[12]) );
  AOI21XL U156 ( .A0(n86), .A1(n67), .B0(n68), .Y(n66) );
  AOI21XL U157 ( .A0(n25), .A1(n170), .B0(n22), .Y(n20) );
  AOI21XL U158 ( .A0(n33), .A1(n171), .B0(n30), .Y(n28) );
  AOI21X1 U159 ( .A0(n45), .A1(n37), .B0(n38), .Y(n36) );
  NOR2XL U160 ( .A(B[5]), .B(A[5]), .Y(n63) );
  NOR2XL U161 ( .A(B[2]), .B(A[2]), .Y(n79) );
  NAND2XL U162 ( .A(B[8]), .B(A[8]), .Y(n51) );
  NOR2X1 U163 ( .A(B[4]), .B(A[4]), .Y(n69) );
  NAND2XL U164 ( .A(B[4]), .B(A[4]), .Y(n70) );
  NAND2XL U165 ( .A(B[6]), .B(A[6]), .Y(n59) );
  NAND2XL U166 ( .A(B[2]), .B(A[2]), .Y(n80) );
  NOR2X1 U167 ( .A(B[1]), .B(A[1]), .Y(n87) );
  NAND2XL U168 ( .A(B[1]), .B(A[1]), .Y(n88) );
  NAND2XL U169 ( .A(B[3]), .B(A[3]), .Y(n77) );
  NAND2BXL U170 ( .AN(n89), .B(n90), .Y(n16) );
  NOR2XL U171 ( .A(B[0]), .B(A[0]), .Y(n89) );
  CLKINVX1 U172 ( .A(n66), .Y(n65) );
  CLKINVX1 U173 ( .A(n86), .Y(n85) );
  NAND2X1 U174 ( .A(n97), .B(n43), .Y(n7) );
  CLKINVX1 U175 ( .A(n42), .Y(n97) );
  NOR2X1 U176 ( .A(n72), .B(n69), .Y(n67) );
  NOR2X1 U177 ( .A(n53), .B(n50), .Y(n48) );
  XNOR2X1 U178 ( .A(n52), .B(n8), .Y(SUM[8]) );
  NAND2X1 U179 ( .A(n98), .B(n51), .Y(n8) );
  OAI21XL U180 ( .A0(n55), .A1(n53), .B0(n54), .Y(n52) );
  CLKINVX1 U181 ( .A(n50), .Y(n98) );
  XNOR2X1 U182 ( .A(n41), .B(n6), .Y(SUM[10]) );
  NAND2X1 U183 ( .A(n96), .B(n40), .Y(n6) );
  OAI21XL U184 ( .A0(n44), .A1(n42), .B0(n43), .Y(n41) );
  NAND2X1 U185 ( .A(n170), .B(n24), .Y(n2) );
  NAND2X1 U186 ( .A(n171), .B(n32), .Y(n4) );
  XNOR2X1 U187 ( .A(n78), .B(n13), .Y(SUM[3]) );
  NAND2X1 U188 ( .A(n169), .B(n77), .Y(n13) );
  OAI21XL U189 ( .A0(n85), .A1(n79), .B0(n80), .Y(n78) );
  XNOR2X1 U190 ( .A(n71), .B(n12), .Y(SUM[4]) );
  NAND2X1 U191 ( .A(n102), .B(n70), .Y(n12) );
  OAI21XL U192 ( .A0(n85), .A1(n72), .B0(n73), .Y(n71) );
  CLKINVX1 U193 ( .A(n69), .Y(n102) );
  XNOR2X1 U194 ( .A(n65), .B(n11), .Y(SUM[5]) );
  NAND2X1 U195 ( .A(n61), .B(n64), .Y(n11) );
  OAI21XL U196 ( .A0(n58), .A1(n64), .B0(n59), .Y(n57) );
  AOI21X1 U197 ( .A0(n169), .A1(n82), .B0(n75), .Y(n73) );
  CLKINVX1 U198 ( .A(n80), .Y(n82) );
  CLKINVX1 U199 ( .A(n77), .Y(n75) );
  OAI21XL U200 ( .A0(n36), .A1(n34), .B0(n35), .Y(n33) );
  NOR2X1 U201 ( .A(n42), .B(n39), .Y(n37) );
  OAI21XL U202 ( .A0(n39), .A1(n43), .B0(n40), .Y(n38) );
  CLKINVX1 U203 ( .A(n32), .Y(n30) );
  CLKINVX1 U204 ( .A(n24), .Y(n22) );
  OAI21XL U205 ( .A0(n50), .A1(n54), .B0(n51), .Y(n49) );
  NOR2X1 U206 ( .A(n63), .B(n58), .Y(n56) );
  NAND2X1 U207 ( .A(n169), .B(n81), .Y(n72) );
  AOI21X1 U208 ( .A0(n65), .A1(n61), .B0(n62), .Y(n60) );
  CLKINVX1 U209 ( .A(n79), .Y(n81) );
  CLKINVX1 U210 ( .A(n63), .Y(n61) );
  CLKINVX1 U211 ( .A(n64), .Y(n62) );
  NOR2X1 U212 ( .A(B[9]), .B(A[9]), .Y(n42) );
  NOR2X1 U213 ( .A(B[10]), .B(A[10]), .Y(n39) );
  NOR2X1 U214 ( .A(B[11]), .B(A[11]), .Y(n34) );
  NAND2X1 U215 ( .A(B[12]), .B(A[12]), .Y(n32) );
  NAND2X1 U216 ( .A(B[14]), .B(A[14]), .Y(n24) );
  NAND2X1 U217 ( .A(B[9]), .B(A[9]), .Y(n43) );
  OR2X1 U218 ( .A(B[14]), .B(A[14]), .Y(n170) );
  NAND2X1 U219 ( .A(B[10]), .B(A[10]), .Y(n40) );
  NAND2X1 U220 ( .A(B[11]), .B(A[11]), .Y(n35) );
  OR2X1 U221 ( .A(B[12]), .B(A[12]), .Y(n171) );
  NOR2X1 U222 ( .A(B[13]), .B(A[13]), .Y(n26) );
  NOR2X1 U223 ( .A(B[15]), .B(A[15]), .Y(n18) );
  NAND2X1 U224 ( .A(B[13]), .B(A[13]), .Y(n27) );
  NAND2X1 U225 ( .A(B[15]), .B(A[15]), .Y(n19) );
  CLKINVX1 U226 ( .A(n16), .Y(SUM[0]) );
endmodule


module datapath_DW01_add_8 ( A, B, CI, SUM, CO );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n20,
         n21, n22, n23, n24, n26, n28, n29, n30, n31, n32, n34, n36, n37, n39,
         n40, n42, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n85,
         n86, n87, n88, n89, n94, n102, n165, n167, n168, n169, n170, n171,
         n172, n173, n174, n175;

  XOR2X1 U11 ( .A(n24), .B(n2), .Y(SUM[14]) );
  XOR2X1 U25 ( .A(n32), .B(n4), .Y(SUM[12]) );
  XOR2X1 U39 ( .A(n40), .B(n6), .Y(SUM[10]) );
  XOR2X1 U63 ( .A(n55), .B(n9), .Y(SUM[7]) );
  XOR2X1 U69 ( .A(n60), .B(n10), .Y(SUM[6]) );
  XOR2X1 U104 ( .A(n85), .B(n14), .Y(SUM[2]) );
  XOR2X1 U114 ( .A(n15), .B(n89), .Y(SUM[1]) );
  OAI21X1 U127 ( .A0(n66), .A1(n46), .B0(n47), .Y(n45) );
  AOI21X1 U128 ( .A0(n86), .A1(n67), .B0(n68), .Y(n66) );
  NAND2XL U129 ( .A(B[2]), .B(A[2]), .Y(n80) );
  NAND2X1 U130 ( .A(n168), .B(n39), .Y(n37) );
  NAND2X1 U131 ( .A(n167), .B(n165), .Y(n168) );
  CLKINVX1 U132 ( .A(n40), .Y(n167) );
  OR2X1 U133 ( .A(B[10]), .B(A[10]), .Y(n165) );
  OAI2BB1X1 U134 ( .A0N(n21), .A1N(n174), .B0(n20), .Y(SUM[16]) );
  NOR2XL U135 ( .A(B[2]), .B(A[2]), .Y(n79) );
  OAI21XL U136 ( .A0(n73), .A1(n69), .B0(n70), .Y(n68) );
  AOI21X1 U137 ( .A0(n29), .A1(n175), .B0(n26), .Y(n24) );
  OAI21XL U138 ( .A0(n58), .A1(n64), .B0(n59), .Y(n57) );
  NOR2XL U139 ( .A(n53), .B(n50), .Y(n48) );
  AOI21X1 U140 ( .A0(n57), .A1(n48), .B0(n49), .Y(n47) );
  XNOR2XL U141 ( .A(n21), .B(n1), .Y(SUM[15]) );
  INVX1 U142 ( .A(n76), .Y(n74) );
  NOR2XL U143 ( .A(B[1]), .B(A[1]), .Y(n87) );
  AOI21XL U144 ( .A0(n65), .A1(n56), .B0(n57), .Y(n55) );
  NAND2XL U145 ( .A(n61), .B(n64), .Y(n11) );
  NAND2BX1 U146 ( .AN(n22), .B(n23), .Y(n2) );
  INVXL U147 ( .A(n64), .Y(n62) );
  XNOR2XL U148 ( .A(n29), .B(n3), .Y(SUM[13]) );
  XNOR2XL U149 ( .A(n45), .B(n7), .Y(SUM[9]) );
  NAND2XL U150 ( .A(n173), .B(n44), .Y(n7) );
  NAND2BXL U151 ( .AN(n53), .B(n54), .Y(n9) );
  NAND2BXL U152 ( .AN(n50), .B(n51), .Y(n8) );
  NAND2XL U153 ( .A(n81), .B(n80), .Y(n14) );
  NAND2X1 U154 ( .A(n169), .B(n170), .Y(n171) );
  NAND2X1 U155 ( .A(n171), .B(n23), .Y(n21) );
  INVXL U156 ( .A(n24), .Y(n169) );
  CLKINVX1 U157 ( .A(n22), .Y(n170) );
  NOR2XL U158 ( .A(B[5]), .B(A[5]), .Y(n63) );
  NOR2X1 U159 ( .A(B[6]), .B(A[6]), .Y(n58) );
  NAND2XL U160 ( .A(B[6]), .B(A[6]), .Y(n59) );
  NAND2XL U161 ( .A(B[8]), .B(A[8]), .Y(n51) );
  NOR2X1 U162 ( .A(B[4]), .B(A[4]), .Y(n69) );
  NAND2XL U163 ( .A(B[9]), .B(A[9]), .Y(n44) );
  NAND2XL U164 ( .A(B[3]), .B(A[3]), .Y(n77) );
  NAND2XL U165 ( .A(B[4]), .B(A[4]), .Y(n70) );
  NAND2X1 U166 ( .A(B[14]), .B(A[14]), .Y(n23) );
  NAND2X1 U167 ( .A(B[10]), .B(A[10]), .Y(n39) );
  XNOR2XL U168 ( .A(n37), .B(n5), .Y(SUM[11]) );
  NOR2XL U169 ( .A(B[14]), .B(A[14]), .Y(n22) );
  NAND2XL U170 ( .A(B[1]), .B(A[1]), .Y(n88) );
  CLKINVX1 U171 ( .A(n66), .Y(n65) );
  CLKINVX1 U172 ( .A(n86), .Y(n85) );
  OAI21XL U173 ( .A0(n87), .A1(n89), .B0(n88), .Y(n86) );
  NOR2X1 U174 ( .A(n72), .B(n69), .Y(n67) );
  XNOR2X1 U175 ( .A(n71), .B(n12), .Y(SUM[4]) );
  NAND2X1 U176 ( .A(n102), .B(n70), .Y(n12) );
  OAI21XL U177 ( .A0(n85), .A1(n72), .B0(n73), .Y(n71) );
  CLKINVX1 U178 ( .A(n69), .Y(n102) );
  XNOR2X1 U179 ( .A(n78), .B(n13), .Y(SUM[3]) );
  NAND2X1 U180 ( .A(n74), .B(n77), .Y(n13) );
  OAI21XL U181 ( .A0(n85), .A1(n79), .B0(n80), .Y(n78) );
  XNOR2X1 U182 ( .A(n65), .B(n11), .Y(SUM[5]) );
  AOI21X1 U183 ( .A0(n74), .A1(n82), .B0(n75), .Y(n73) );
  CLKINVX1 U184 ( .A(n77), .Y(n75) );
  CLKINVX1 U185 ( .A(n80), .Y(n82) );
  NAND2X1 U186 ( .A(n56), .B(n48), .Y(n46) );
  OAI21XL U187 ( .A0(n32), .A1(n30), .B0(n31), .Y(n29) );
  AOI21X1 U188 ( .A0(n45), .A1(n173), .B0(n42), .Y(n40) );
  CLKINVX1 U189 ( .A(n44), .Y(n42) );
  AOI21X1 U190 ( .A0(n37), .A1(n172), .B0(n34), .Y(n32) );
  CLKINVX1 U191 ( .A(n36), .Y(n34) );
  CLKINVX1 U192 ( .A(n28), .Y(n26) );
  OAI21XL U193 ( .A0(n50), .A1(n54), .B0(n51), .Y(n49) );
  NOR2X1 U194 ( .A(n63), .B(n58), .Y(n56) );
  OAI21XL U195 ( .A0(n55), .A1(n53), .B0(n54), .Y(n52) );
  NAND2X1 U196 ( .A(n74), .B(n81), .Y(n72) );
  AOI21X1 U197 ( .A0(n65), .A1(n61), .B0(n62), .Y(n60) );
  CLKINVX1 U198 ( .A(n79), .Y(n81) );
  NAND2X1 U199 ( .A(n175), .B(n28), .Y(n3) );
  NAND2X1 U200 ( .A(n172), .B(n36), .Y(n5) );
  NAND2X1 U201 ( .A(n174), .B(n20), .Y(n1) );
  NAND2BX1 U202 ( .AN(n87), .B(n88), .Y(n15) );
  CLKINVX1 U203 ( .A(n30), .Y(n94) );
  CLKINVX1 U204 ( .A(n63), .Y(n61) );
  NAND2BX1 U205 ( .AN(n58), .B(n59), .Y(n10) );
  NOR2X1 U206 ( .A(B[7]), .B(A[7]), .Y(n53) );
  NOR2X1 U207 ( .A(B[0]), .B(A[0]), .Y(n89) );
  NOR2X1 U208 ( .A(B[8]), .B(A[8]), .Y(n50) );
  NOR2X1 U209 ( .A(B[12]), .B(A[12]), .Y(n30) );
  XNOR2X1 U210 ( .A(n52), .B(n8), .Y(SUM[8]) );
  NAND2X1 U211 ( .A(B[5]), .B(A[5]), .Y(n64) );
  NAND2X1 U212 ( .A(B[7]), .B(A[7]), .Y(n54) );
  NAND2X1 U213 ( .A(B[12]), .B(A[12]), .Y(n31) );
  NAND2X1 U214 ( .A(B[11]), .B(A[11]), .Y(n36) );
  NAND2X1 U215 ( .A(n94), .B(n31), .Y(n4) );
  NAND2X1 U216 ( .A(n165), .B(n39), .Y(n6) );
  NOR2X1 U217 ( .A(B[3]), .B(A[3]), .Y(n76) );
  OR2X1 U218 ( .A(B[11]), .B(A[11]), .Y(n172) );
  OR2X1 U219 ( .A(B[9]), .B(A[9]), .Y(n173) );
  NAND2X1 U220 ( .A(B[15]), .B(A[15]), .Y(n20) );
  NAND2X1 U221 ( .A(B[13]), .B(A[13]), .Y(n28) );
  OR2X1 U222 ( .A(B[15]), .B(A[15]), .Y(n174) );
  OR2X1 U223 ( .A(B[13]), .B(A[13]), .Y(n175) );
  XNOR2XL U224 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module datapath_DW01_add_7 ( A, B, CI, SUM, CO );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n21, n22, n23, n24, n25, n27, n29, n30, n31, n32, n33, n35, n37, n38,
         n39, n40, n41, n43, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n76, n78, n79, n80, n81, n82, n83, n86,
         n87, n88, n89, n90, n91, n96, n98, n101, n102, n107, n168, n169, n170,
         n171, n172;

  XOR2X1 U11 ( .A(n25), .B(n2), .Y(SUM[14]) );
  XOR2X1 U25 ( .A(n33), .B(n4), .Y(SUM[12]) );
  XOR2X1 U39 ( .A(n41), .B(n6), .Y(SUM[10]) );
  XOR2X1 U63 ( .A(n56), .B(n9), .Y(SUM[7]) );
  XOR2X1 U69 ( .A(n61), .B(n10), .Y(SUM[6]) );
  XOR2X1 U104 ( .A(n86), .B(n14), .Y(SUM[2]) );
  XOR2X1 U114 ( .A(n15), .B(n91), .Y(SUM[1]) );
  AOI21XL U129 ( .A0(n46), .A1(n170), .B0(n43), .Y(n41) );
  OAI21XL U130 ( .A0(n67), .A1(n47), .B0(n48), .Y(n46) );
  OAI21XL U131 ( .A0(n25), .A1(n23), .B0(n24), .Y(n22) );
  OAI2BB1XL U132 ( .A0N(n22), .A1N(n172), .B0(n21), .Y(SUM[16]) );
  OAI21XL U133 ( .A0(n88), .A1(n91), .B0(n89), .Y(n87) );
  OR2X1 U134 ( .A(B[3]), .B(A[3]), .Y(n168) );
  AOI21XL U135 ( .A0(n58), .A1(n49), .B0(n50), .Y(n48) );
  INVXL U136 ( .A(n87), .Y(n86) );
  AOI21XL U137 ( .A0(n87), .A1(n68), .B0(n69), .Y(n67) );
  OAI21X2 U138 ( .A0(n33), .A1(n31), .B0(n32), .Y(n30) );
  AOI21X1 U139 ( .A0(n38), .A1(n169), .B0(n35), .Y(n33) );
  OAI21XL U140 ( .A0(n74), .A1(n70), .B0(n71), .Y(n69) );
  XNOR2X1 U141 ( .A(n30), .B(n3), .Y(SUM[13]) );
  NAND2BXL U142 ( .AN(n90), .B(n91), .Y(n16) );
  AOI21X1 U143 ( .A0(n30), .A1(n171), .B0(n27), .Y(n25) );
  NOR2X1 U144 ( .A(B[4]), .B(A[4]), .Y(n70) );
  NAND2X1 U145 ( .A(B[5]), .B(A[5]), .Y(n65) );
  AOI21XL U146 ( .A0(n66), .A1(n57), .B0(n58), .Y(n56) );
  NAND2BX1 U147 ( .AN(n23), .B(n24), .Y(n2) );
  NAND2XL U148 ( .A(n82), .B(n81), .Y(n14) );
  XNOR2XL U149 ( .A(n38), .B(n5), .Y(SUM[11]) );
  XNOR2XL U150 ( .A(n46), .B(n7), .Y(SUM[9]) );
  NOR2XL U151 ( .A(B[7]), .B(A[7]), .Y(n54) );
  NOR2XL U152 ( .A(B[8]), .B(A[8]), .Y(n51) );
  NOR2XL U153 ( .A(B[5]), .B(A[5]), .Y(n64) );
  NOR2XL U154 ( .A(B[2]), .B(A[2]), .Y(n80) );
  NOR2X1 U155 ( .A(B[6]), .B(A[6]), .Y(n59) );
  NAND2XL U156 ( .A(B[0]), .B(A[0]), .Y(n91) );
  NAND2XL U157 ( .A(B[7]), .B(A[7]), .Y(n55) );
  NAND2XL U158 ( .A(B[6]), .B(A[6]), .Y(n60) );
  NAND2XL U159 ( .A(B[8]), .B(A[8]), .Y(n52) );
  NAND2XL U160 ( .A(B[9]), .B(A[9]), .Y(n45) );
  NAND2XL U161 ( .A(B[3]), .B(A[3]), .Y(n78) );
  NAND2XL U162 ( .A(B[2]), .B(A[2]), .Y(n81) );
  NAND2XL U163 ( .A(B[4]), .B(A[4]), .Y(n71) );
  OR2XL U164 ( .A(B[9]), .B(A[9]), .Y(n170) );
  NOR2XL U165 ( .A(B[0]), .B(A[0]), .Y(n90) );
  NAND2XL U166 ( .A(B[1]), .B(A[1]), .Y(n89) );
  NOR2XL U167 ( .A(B[1]), .B(A[1]), .Y(n88) );
  OAI21XL U168 ( .A0(n86), .A1(n73), .B0(n74), .Y(n72) );
  CLKINVX1 U169 ( .A(n67), .Y(n66) );
  NOR2X1 U170 ( .A(n73), .B(n70), .Y(n68) );
  NAND2X1 U171 ( .A(n102), .B(n60), .Y(n10) );
  OAI21XL U172 ( .A0(n59), .A1(n65), .B0(n60), .Y(n58) );
  AOI21X1 U173 ( .A0(n168), .A1(n83), .B0(n76), .Y(n74) );
  CLKINVX1 U174 ( .A(n78), .Y(n76) );
  CLKINVX1 U175 ( .A(n81), .Y(n83) );
  NAND2X1 U176 ( .A(n57), .B(n49), .Y(n47) );
  NOR2X1 U177 ( .A(n54), .B(n51), .Y(n49) );
  OAI21XL U178 ( .A0(n41), .A1(n39), .B0(n40), .Y(n38) );
  CLKINVX1 U179 ( .A(n45), .Y(n43) );
  CLKINVX1 U180 ( .A(n37), .Y(n35) );
  CLKINVX1 U181 ( .A(n29), .Y(n27) );
  OAI21XL U182 ( .A0(n51), .A1(n55), .B0(n52), .Y(n50) );
  NOR2X1 U183 ( .A(n64), .B(n59), .Y(n57) );
  OAI21XL U184 ( .A0(n56), .A1(n54), .B0(n55), .Y(n53) );
  OAI21XL U185 ( .A0(n86), .A1(n80), .B0(n81), .Y(n79) );
  NAND2X1 U186 ( .A(n168), .B(n82), .Y(n73) );
  AOI21X1 U187 ( .A0(n66), .A1(n62), .B0(n63), .Y(n61) );
  CLKINVX1 U188 ( .A(n65), .Y(n63) );
  NAND2X1 U189 ( .A(n96), .B(n32), .Y(n4) );
  NAND2X1 U190 ( .A(n101), .B(n55), .Y(n9) );
  NAND2X1 U191 ( .A(n98), .B(n40), .Y(n6) );
  XNOR2X1 U192 ( .A(n53), .B(n8), .Y(SUM[8]) );
  XNOR2X1 U193 ( .A(n79), .B(n13), .Y(SUM[3]) );
  XNOR2X1 U194 ( .A(n72), .B(n12), .Y(SUM[4]) );
  XNOR2X1 U195 ( .A(n66), .B(n11), .Y(SUM[5]) );
  CLKINVX1 U196 ( .A(n80), .Y(n82) );
  CLKINVX1 U197 ( .A(n88), .Y(n107) );
  NAND2X1 U198 ( .A(n107), .B(n89), .Y(n15) );
  CLKINVX1 U199 ( .A(n31), .Y(n96) );
  NAND2X1 U200 ( .A(n169), .B(n37), .Y(n5) );
  NAND2X1 U201 ( .A(n170), .B(n45), .Y(n7) );
  NAND2X1 U202 ( .A(n171), .B(n29), .Y(n3) );
  XNOR2X1 U203 ( .A(n22), .B(n1), .Y(SUM[15]) );
  NAND2X1 U204 ( .A(n172), .B(n21), .Y(n1) );
  NAND2X1 U205 ( .A(n62), .B(n65), .Y(n11) );
  CLKINVX1 U206 ( .A(n16), .Y(SUM[0]) );
  CLKINVX1 U207 ( .A(n64), .Y(n62) );
  NAND2X1 U208 ( .A(n168), .B(n78), .Y(n13) );
  CLKINVX1 U209 ( .A(n54), .Y(n101) );
  NAND2BX1 U210 ( .AN(n70), .B(n71), .Y(n12) );
  CLKINVX1 U211 ( .A(n59), .Y(n102) );
  NAND2BX1 U212 ( .AN(n51), .B(n52), .Y(n8) );
  CLKINVX1 U213 ( .A(n39), .Y(n98) );
  NOR2X1 U214 ( .A(B[12]), .B(A[12]), .Y(n31) );
  NOR2X1 U215 ( .A(B[10]), .B(A[10]), .Y(n39) );
  NAND2X1 U216 ( .A(B[12]), .B(A[12]), .Y(n32) );
  NAND2X1 U217 ( .A(B[11]), .B(A[11]), .Y(n37) );
  NAND2X1 U218 ( .A(B[10]), .B(A[10]), .Y(n40) );
  OR2X1 U219 ( .A(B[11]), .B(A[11]), .Y(n169) );
  NOR2X1 U220 ( .A(B[14]), .B(A[14]), .Y(n23) );
  NAND2X1 U221 ( .A(B[15]), .B(A[15]), .Y(n21) );
  OR2X1 U222 ( .A(B[13]), .B(A[13]), .Y(n171) );
  NAND2X1 U223 ( .A(B[13]), .B(A[13]), .Y(n29) );
  NAND2X1 U224 ( .A(B[14]), .B(A[14]), .Y(n24) );
  OR2X1 U225 ( .A(B[15]), .B(A[15]), .Y(n172) );
endmodule


module datapath ( V, C, N, Z, R0, R1, R2, R3, R4, R5, R6, R7, R8, R9, R10, R11, 
        R12, R13, R14, R15, BUSA, BUSB, control, constant, data, clk, rst_n );
  output [15:0] R0;
  output [15:0] R1;
  output [15:0] R2;
  output [15:0] R3;
  output [15:0] R4;
  output [15:0] R5;
  output [15:0] R6;
  output [15:0] R7;
  output [15:0] R8;
  output [15:0] R9;
  output [15:0] R10;
  output [15:0] R11;
  output [15:0] R12;
  output [15:0] R13;
  output [15:0] R14;
  output [15:0] R15;
  output [15:0] BUSA;
  output [15:0] BUSB;
  input [25:0] control;
  input [15:0] constant;
  input [15:0] data;
  input clk, rst_n;
  output V, C, N, Z;
  wire   N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, N67, N68, N69,
         N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N101,
         N102, N103, N104, N105, N106, N107, N109, N110, N111, N112, N113,
         N114, N115, \FUResult[15] , N201, N202, N203, N204, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N294, N295, N296, N297, N298, N299, N300, N301, N302,
         N303, N304, N305, N306, N307, N308, N309, N433, N434, N435, N436,
         N437, N438, N439, N440, N441, N442, N443, N444, N445, N446, N447,
         N448, N449, N452, N453, N454, N455, N456, N457, N458, N459, N460,
         N461, N462, N463, N464, N465, N466, N467, N468, N491, N492, N493,
         N494, N495, N496, N497, N498, N499, N500, N501, N502, N503, N504,
         N505, N506, N507, N513, N514, N515, N516, N517, N518, N519, N520,
         N521, N522, N523, N524, N525, N526, N527, N528, N529, N552, N553,
         N554, N555, N556, N557, N558, N559, N560, N561, N562, N563, N564,
         N565, N566, N567, N568, n41, n47, n48, n49, n50, n51, n52, n53, n54,
         n69, n71, n72, n73, n74, n75, n76, n77, n78, n85, n86, n87, n88, n90,
         n91, n93, n94, n95, n97, n98, n100, n103, n105, n106, n108, n110,
         n112, n113, n115, n118, n121, n123, n126, n128, n129, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, \add_233/carry[2] , \add_233/carry[3] ,
         \add_233/carry[4] , \add_233/carry[5] , \add_233/carry[6] ,
         \add_233/carry[7] , \add_233/carry[8] , n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868;
  wire   [15:0] MUXB;
  assign N53 = control[22];
  assign N54 = control[23];
  assign N55 = control[24];
  assign N56 = control[25];
  assign N57 = control[14];
  assign N58 = control[15];
  assign N59 = control[16];
  assign N60 = control[17];
  assign N61 = control[18];
  assign N62 = control[19];
  assign N63 = control[20];
  assign N64 = control[21];
  assign N = \FUResult[15] ;
  assign N201 = control[2];

  datapath_DW01_inc_0 add_170 ( .A({1'b0, BUSA}), .SUM({N449, N448, N447, N446, 
        N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, 
        N433}) );
  datapath_DW_rightsh_1 srl_143 ( .A({n870, MUXB[14:12], n852, MUXB[10:1], 
        n851}), .DATA_TC(1'b0), .SH({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n1865, N204, N203, 
        N202, N201}), .B({N309, N308, N307, N306, N305, N304, N303, N302, N301, 
        N300, N299, N298, N297, N296, N295, N294}) );
  datapath_DW_leftsh_0 sll_133 ( .A({n870, MUXB[14:12], n852, MUXB[10:1], n851}), .SH({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, n1865, N204, N203, N202, N201}), .B({N222, N221, 
        N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, 
        N208, N207}) );
  datapath_DW01_add_5 add_1_root_add_220_2 ( .A({1'b0, BUSA}), .B({1'b0, n891, 
        n886, n890, n882, n885, n884, n888, n883, n887, n878, n879, n881, n876, 
        n877, n880, n889}), .CI(1'b1), .SUM({N568, N567, N566, N565, N564, 
        N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552}) );
  datapath_DW01_add_6 add_206 ( .A({1'b0, BUSA}), .B({1'b0, n891, n886, n890, 
        n882, n885, n884, n888, n883, n887, n878, n879, n881, n876, n877, n880, 
        n889}), .CI(1'b0), .SUM({N529, N528, N527, N526, N525, N524, N523, 
        N522, N521, N520, N519, N518, N517, N516, N515, N514, N513}) );
  datapath_DW01_add_8 add_1_root_add_192_2 ( .A({1'b0, BUSA}), .B({1'b0, BUSB}), .CI(1'b1), .SUM({N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, 
        N497, N496, N495, N494, N493, N492, N491}) );
  datapath_DW01_add_7 add_179 ( .A({1'b0, BUSA}), .B({1'b0, BUSB}), .CI(1'b0), 
        .SUM({N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, 
        N457, N456, N455, N454, N453, N452}) );
  DFFRX1 \R_reg[3][15]  ( .D(n787), .CK(clk), .RN(rst_n), .Q(R3[15]), .QN(n531) );
  DFFRX1 \R_reg[3][14]  ( .D(n786), .CK(clk), .RN(rst_n), .Q(R3[14]), .QN(n530) );
  DFFRX1 \R_reg[3][13]  ( .D(n785), .CK(clk), .RN(rst_n), .Q(R3[13]), .QN(n529) );
  DFFRX1 \R_reg[3][12]  ( .D(n784), .CK(clk), .RN(rst_n), .Q(R3[12]), .QN(n528) );
  DFFRX1 \R_reg[3][11]  ( .D(n783), .CK(clk), .RN(rst_n), .Q(R3[11]), .QN(n527) );
  DFFRX1 \R_reg[3][10]  ( .D(n782), .CK(clk), .RN(rst_n), .Q(R3[10]), .QN(n526) );
  DFFRX1 \R_reg[3][9]  ( .D(n781), .CK(clk), .RN(rst_n), .Q(R3[9]), .QN(n525)
         );
  DFFRX1 \R_reg[3][6]  ( .D(n778), .CK(clk), .RN(rst_n), .Q(R3[6]), .QN(n522)
         );
  DFFRX1 \R_reg[3][5]  ( .D(n777), .CK(clk), .RN(rst_n), .Q(R3[5]), .QN(n521)
         );
  DFFRX1 \R_reg[3][0]  ( .D(n772), .CK(clk), .RN(rst_n), .Q(R3[0]), .QN(n516)
         );
  DFFRX1 \R_reg[7][15]  ( .D(n723), .CK(clk), .RN(rst_n), .Q(R7[15]), .QN(n467) );
  DFFRX1 \R_reg[7][14]  ( .D(n722), .CK(clk), .RN(rst_n), .Q(R7[14]), .QN(n466) );
  DFFRX1 \R_reg[7][13]  ( .D(n721), .CK(clk), .RN(rst_n), .Q(R7[13]), .QN(n465) );
  DFFRX1 \R_reg[7][12]  ( .D(n720), .CK(clk), .RN(rst_n), .Q(R7[12]), .QN(n464) );
  DFFRX1 \R_reg[7][11]  ( .D(n719), .CK(clk), .RN(rst_n), .Q(R7[11]), .QN(n463) );
  DFFRX1 \R_reg[7][10]  ( .D(n718), .CK(clk), .RN(rst_n), .Q(R7[10]), .QN(n462) );
  DFFRX1 \R_reg[7][9]  ( .D(n717), .CK(clk), .RN(rst_n), .Q(R7[9]), .QN(n461)
         );
  DFFRX1 \R_reg[7][8]  ( .D(n716), .CK(clk), .RN(rst_n), .Q(R7[8]), .QN(n460)
         );
  DFFRX1 \R_reg[7][7]  ( .D(n715), .CK(clk), .RN(rst_n), .Q(R7[7]), .QN(n459)
         );
  DFFRX1 \R_reg[7][6]  ( .D(n714), .CK(clk), .RN(rst_n), .Q(R7[6]), .QN(n458)
         );
  DFFRX1 \R_reg[7][5]  ( .D(n713), .CK(clk), .RN(rst_n), .Q(R7[5]), .QN(n457)
         );
  DFFRX1 \R_reg[7][0]  ( .D(n708), .CK(clk), .RN(rst_n), .Q(R7[0]), .QN(n452)
         );
  DFFRX1 \R_reg[11][15]  ( .D(n659), .CK(clk), .RN(rst_n), .Q(R11[15]), .QN(
        n403) );
  DFFRX1 \R_reg[11][14]  ( .D(n658), .CK(clk), .RN(rst_n), .Q(R11[14]), .QN(
        n402) );
  DFFRX1 \R_reg[11][13]  ( .D(n657), .CK(clk), .RN(rst_n), .Q(R11[13]), .QN(
        n401) );
  DFFRX1 \R_reg[11][12]  ( .D(n656), .CK(clk), .RN(rst_n), .Q(R11[12]), .QN(
        n400) );
  DFFRX1 \R_reg[11][11]  ( .D(n655), .CK(clk), .RN(rst_n), .Q(R11[11]), .QN(
        n399) );
  DFFRX1 \R_reg[11][10]  ( .D(n654), .CK(clk), .RN(rst_n), .Q(R11[10]), .QN(
        n398) );
  DFFRX1 \R_reg[11][9]  ( .D(n653), .CK(clk), .RN(rst_n), .Q(R11[9]), .QN(n397) );
  DFFRX1 \R_reg[11][6]  ( .D(n650), .CK(clk), .RN(rst_n), .Q(R11[6]), .QN(n394) );
  DFFRX1 \R_reg[11][5]  ( .D(n649), .CK(clk), .RN(rst_n), .Q(R11[5]), .QN(n393) );
  DFFRX1 \R_reg[11][0]  ( .D(n644), .CK(clk), .RN(rst_n), .Q(R11[0]), .QN(n388) );
  DFFRX1 \R_reg[15][15]  ( .D(n595), .CK(clk), .RN(rst_n), .Q(R15[15]), .QN(
        n339) );
  DFFRX1 \R_reg[15][14]  ( .D(n594), .CK(clk), .RN(rst_n), .Q(R15[14]), .QN(
        n338) );
  DFFRX1 \R_reg[15][13]  ( .D(n593), .CK(clk), .RN(rst_n), .Q(R15[13]), .QN(
        n337) );
  DFFRX1 \R_reg[15][12]  ( .D(n592), .CK(clk), .RN(rst_n), .Q(R15[12]), .QN(
        n336) );
  DFFRX1 \R_reg[15][11]  ( .D(n591), .CK(clk), .RN(rst_n), .Q(R15[11]), .QN(
        n335) );
  DFFRX1 \R_reg[15][10]  ( .D(n590), .CK(clk), .RN(rst_n), .Q(R15[10]), .QN(
        n334) );
  DFFRX1 \R_reg[15][9]  ( .D(n589), .CK(clk), .RN(rst_n), .Q(R15[9]), .QN(n333) );
  DFFRX1 \R_reg[15][8]  ( .D(n588), .CK(clk), .RN(rst_n), .Q(R15[8]), .QN(n332) );
  DFFRX1 \R_reg[15][7]  ( .D(n587), .CK(clk), .RN(rst_n), .Q(R15[7]), .QN(n331) );
  DFFRX1 \R_reg[15][6]  ( .D(n586), .CK(clk), .RN(rst_n), .Q(R15[6]), .QN(n330) );
  DFFRX1 \R_reg[15][5]  ( .D(n585), .CK(clk), .RN(rst_n), .Q(R15[5]), .QN(n329) );
  DFFRX1 \R_reg[15][0]  ( .D(n580), .CK(clk), .RN(rst_n), .Q(R15[0]), .QN(n324) );
  DFFRX1 \R_reg[1][15]  ( .D(n819), .CK(clk), .RN(rst_n), .Q(R1[15]), .QN(n563) );
  DFFRX1 \R_reg[1][14]  ( .D(n818), .CK(clk), .RN(rst_n), .Q(R1[14]), .QN(n562) );
  DFFRX1 \R_reg[1][13]  ( .D(n817), .CK(clk), .RN(rst_n), .Q(R1[13]), .QN(n561) );
  DFFRX1 \R_reg[1][12]  ( .D(n816), .CK(clk), .RN(rst_n), .Q(R1[12]), .QN(n560) );
  DFFRX1 \R_reg[1][11]  ( .D(n815), .CK(clk), .RN(rst_n), .Q(R1[11]), .QN(n559) );
  DFFRX1 \R_reg[1][10]  ( .D(n814), .CK(clk), .RN(rst_n), .Q(R1[10]), .QN(n558) );
  DFFRX1 \R_reg[1][9]  ( .D(n813), .CK(clk), .RN(rst_n), .Q(R1[9]), .QN(n557)
         );
  DFFRX1 \R_reg[1][6]  ( .D(n810), .CK(clk), .RN(rst_n), .Q(R1[6]), .QN(n554)
         );
  DFFRX1 \R_reg[1][5]  ( .D(n809), .CK(clk), .RN(rst_n), .Q(R1[5]), .QN(n553)
         );
  DFFRX1 \R_reg[1][0]  ( .D(n804), .CK(clk), .RN(rst_n), .Q(R1[0]), .QN(n548)
         );
  DFFRX1 \R_reg[5][15]  ( .D(n755), .CK(clk), .RN(rst_n), .Q(R5[15]), .QN(n499) );
  DFFRX1 \R_reg[5][14]  ( .D(n754), .CK(clk), .RN(rst_n), .Q(R5[14]), .QN(n498) );
  DFFRX1 \R_reg[5][13]  ( .D(n753), .CK(clk), .RN(rst_n), .Q(R5[13]), .QN(n497) );
  DFFRX1 \R_reg[5][12]  ( .D(n752), .CK(clk), .RN(rst_n), .Q(R5[12]), .QN(n496) );
  DFFRX1 \R_reg[5][11]  ( .D(n751), .CK(clk), .RN(rst_n), .Q(R5[11]), .QN(n495) );
  DFFRX1 \R_reg[5][10]  ( .D(n750), .CK(clk), .RN(rst_n), .Q(R5[10]), .QN(n494) );
  DFFRX1 \R_reg[5][9]  ( .D(n749), .CK(clk), .RN(rst_n), .Q(R5[9]), .QN(n493)
         );
  DFFRX1 \R_reg[5][6]  ( .D(n746), .CK(clk), .RN(rst_n), .Q(R5[6]), .QN(n490)
         );
  DFFRX1 \R_reg[5][5]  ( .D(n745), .CK(clk), .RN(rst_n), .Q(R5[5]), .QN(n489)
         );
  DFFRX1 \R_reg[5][0]  ( .D(n740), .CK(clk), .RN(rst_n), .Q(R5[0]), .QN(n484)
         );
  DFFRX1 \R_reg[9][15]  ( .D(n691), .CK(clk), .RN(rst_n), .Q(R9[15]), .QN(n435) );
  DFFRX1 \R_reg[9][14]  ( .D(n690), .CK(clk), .RN(rst_n), .Q(R9[14]), .QN(n434) );
  DFFRX1 \R_reg[9][13]  ( .D(n689), .CK(clk), .RN(rst_n), .Q(R9[13]), .QN(n433) );
  DFFRX1 \R_reg[9][12]  ( .D(n688), .CK(clk), .RN(rst_n), .Q(R9[12]), .QN(n432) );
  DFFRX1 \R_reg[9][11]  ( .D(n687), .CK(clk), .RN(rst_n), .Q(R9[11]), .QN(n431) );
  DFFRX1 \R_reg[9][10]  ( .D(n686), .CK(clk), .RN(rst_n), .Q(R9[10]), .QN(n430) );
  DFFRX1 \R_reg[9][9]  ( .D(n685), .CK(clk), .RN(rst_n), .Q(R9[9]), .QN(n429)
         );
  DFFRX1 \R_reg[9][6]  ( .D(n682), .CK(clk), .RN(rst_n), .Q(R9[6]), .QN(n426)
         );
  DFFRX1 \R_reg[9][5]  ( .D(n681), .CK(clk), .RN(rst_n), .Q(R9[5]), .QN(n425)
         );
  DFFRX1 \R_reg[9][0]  ( .D(n676), .CK(clk), .RN(rst_n), .Q(R9[0]), .QN(n420)
         );
  DFFRX1 \R_reg[13][15]  ( .D(n627), .CK(clk), .RN(rst_n), .Q(R13[15]), .QN(
        n371) );
  DFFRX1 \R_reg[13][14]  ( .D(n626), .CK(clk), .RN(rst_n), .Q(R13[14]), .QN(
        n370) );
  DFFRX1 \R_reg[13][13]  ( .D(n625), .CK(clk), .RN(rst_n), .Q(R13[13]), .QN(
        n369) );
  DFFRX1 \R_reg[13][12]  ( .D(n624), .CK(clk), .RN(rst_n), .Q(R13[12]), .QN(
        n368) );
  DFFRX1 \R_reg[13][11]  ( .D(n623), .CK(clk), .RN(rst_n), .Q(R13[11]), .QN(
        n367) );
  DFFRX1 \R_reg[13][10]  ( .D(n622), .CK(clk), .RN(rst_n), .Q(R13[10]), .QN(
        n366) );
  DFFRX1 \R_reg[13][9]  ( .D(n621), .CK(clk), .RN(rst_n), .Q(R13[9]), .QN(n365) );
  DFFRX1 \R_reg[13][6]  ( .D(n618), .CK(clk), .RN(rst_n), .Q(R13[6]), .QN(n362) );
  DFFRX1 \R_reg[13][5]  ( .D(n617), .CK(clk), .RN(rst_n), .Q(R13[5]), .QN(n361) );
  DFFRX1 \R_reg[13][0]  ( .D(n612), .CK(clk), .RN(rst_n), .Q(R13[0]), .QN(n356) );
  DFFRX1 \R_reg[0][15]  ( .D(n835), .CK(clk), .RN(rst_n), .Q(R0[15]), .QN(n579) );
  DFFRX1 \R_reg[0][14]  ( .D(n834), .CK(clk), .RN(rst_n), .Q(R0[14]), .QN(n578) );
  DFFRX1 \R_reg[0][13]  ( .D(n833), .CK(clk), .RN(rst_n), .Q(R0[13]), .QN(n577) );
  DFFRX1 \R_reg[0][12]  ( .D(n832), .CK(clk), .RN(rst_n), .Q(R0[12]), .QN(n576) );
  DFFRX1 \R_reg[0][11]  ( .D(n831), .CK(clk), .RN(rst_n), .Q(R0[11]), .QN(n575) );
  DFFRX1 \R_reg[0][10]  ( .D(n830), .CK(clk), .RN(rst_n), .Q(R0[10]), .QN(n574) );
  DFFRX1 \R_reg[0][9]  ( .D(n829), .CK(clk), .RN(rst_n), .Q(R0[9]), .QN(n573)
         );
  DFFRX1 \R_reg[0][6]  ( .D(n826), .CK(clk), .RN(rst_n), .Q(R0[6]), .QN(n570)
         );
  DFFRX1 \R_reg[0][5]  ( .D(n825), .CK(clk), .RN(rst_n), .Q(R0[5]), .QN(n569)
         );
  DFFRX1 \R_reg[0][0]  ( .D(n820), .CK(clk), .RN(rst_n), .Q(R0[0]), .QN(n564)
         );
  DFFRX1 \R_reg[4][15]  ( .D(n771), .CK(clk), .RN(rst_n), .Q(R4[15]), .QN(n515) );
  DFFRX1 \R_reg[4][14]  ( .D(n770), .CK(clk), .RN(rst_n), .Q(R4[14]), .QN(n514) );
  DFFRX1 \R_reg[4][13]  ( .D(n769), .CK(clk), .RN(rst_n), .Q(R4[13]), .QN(n513) );
  DFFRX1 \R_reg[4][12]  ( .D(n768), .CK(clk), .RN(rst_n), .Q(R4[12]), .QN(n512) );
  DFFRX1 \R_reg[4][11]  ( .D(n767), .CK(clk), .RN(rst_n), .Q(R4[11]), .QN(n511) );
  DFFRX1 \R_reg[4][10]  ( .D(n766), .CK(clk), .RN(rst_n), .Q(R4[10]), .QN(n510) );
  DFFRX1 \R_reg[4][9]  ( .D(n765), .CK(clk), .RN(rst_n), .Q(R4[9]), .QN(n509)
         );
  DFFRX1 \R_reg[4][6]  ( .D(n762), .CK(clk), .RN(rst_n), .Q(R4[6]), .QN(n506)
         );
  DFFRX1 \R_reg[4][5]  ( .D(n761), .CK(clk), .RN(rst_n), .Q(R4[5]), .QN(n505)
         );
  DFFRX1 \R_reg[4][0]  ( .D(n756), .CK(clk), .RN(rst_n), .Q(R4[0]), .QN(n500)
         );
  DFFRX1 \R_reg[8][15]  ( .D(n707), .CK(clk), .RN(rst_n), .Q(R8[15]), .QN(n451) );
  DFFRX1 \R_reg[8][14]  ( .D(n706), .CK(clk), .RN(rst_n), .Q(R8[14]), .QN(n450) );
  DFFRX1 \R_reg[8][13]  ( .D(n705), .CK(clk), .RN(rst_n), .Q(R8[13]), .QN(n449) );
  DFFRX1 \R_reg[8][12]  ( .D(n704), .CK(clk), .RN(rst_n), .Q(R8[12]), .QN(n448) );
  DFFRX1 \R_reg[8][11]  ( .D(n703), .CK(clk), .RN(rst_n), .Q(R8[11]), .QN(n447) );
  DFFRX1 \R_reg[8][10]  ( .D(n702), .CK(clk), .RN(rst_n), .Q(R8[10]), .QN(n446) );
  DFFRX1 \R_reg[8][9]  ( .D(n701), .CK(clk), .RN(rst_n), .Q(R8[9]), .QN(n445)
         );
  DFFRX1 \R_reg[8][6]  ( .D(n698), .CK(clk), .RN(rst_n), .Q(R8[6]), .QN(n442)
         );
  DFFRX1 \R_reg[8][5]  ( .D(n697), .CK(clk), .RN(rst_n), .Q(R8[5]), .QN(n441)
         );
  DFFRX1 \R_reg[8][0]  ( .D(n692), .CK(clk), .RN(rst_n), .Q(R8[0]), .QN(n436)
         );
  DFFRX1 \R_reg[12][15]  ( .D(n643), .CK(clk), .RN(rst_n), .Q(R12[15]), .QN(
        n387) );
  DFFRX1 \R_reg[12][14]  ( .D(n642), .CK(clk), .RN(rst_n), .Q(R12[14]), .QN(
        n386) );
  DFFRX1 \R_reg[12][13]  ( .D(n641), .CK(clk), .RN(rst_n), .Q(R12[13]), .QN(
        n385) );
  DFFRX1 \R_reg[12][12]  ( .D(n640), .CK(clk), .RN(rst_n), .Q(R12[12]), .QN(
        n384) );
  DFFRX1 \R_reg[12][11]  ( .D(n639), .CK(clk), .RN(rst_n), .Q(R12[11]), .QN(
        n383) );
  DFFRX1 \R_reg[12][10]  ( .D(n638), .CK(clk), .RN(rst_n), .Q(R12[10]), .QN(
        n382) );
  DFFRX1 \R_reg[12][9]  ( .D(n637), .CK(clk), .RN(rst_n), .Q(R12[9]), .QN(n381) );
  DFFRX1 \R_reg[12][6]  ( .D(n634), .CK(clk), .RN(rst_n), .Q(R12[6]), .QN(n378) );
  DFFRX1 \R_reg[12][5]  ( .D(n633), .CK(clk), .RN(rst_n), .Q(R12[5]), .QN(n377) );
  DFFRX1 \R_reg[12][0]  ( .D(n628), .CK(clk), .RN(rst_n), .Q(R12[0]), .QN(n372) );
  DFFRX1 \R_reg[2][15]  ( .D(n803), .CK(clk), .RN(rst_n), .Q(R2[15]), .QN(n547) );
  DFFRX1 \R_reg[2][14]  ( .D(n802), .CK(clk), .RN(rst_n), .Q(R2[14]), .QN(n546) );
  DFFRX1 \R_reg[2][13]  ( .D(n801), .CK(clk), .RN(rst_n), .Q(R2[13]), .QN(n545) );
  DFFRX1 \R_reg[2][12]  ( .D(n800), .CK(clk), .RN(rst_n), .Q(R2[12]), .QN(n544) );
  DFFRX1 \R_reg[2][11]  ( .D(n799), .CK(clk), .RN(rst_n), .Q(R2[11]), .QN(n543) );
  DFFRX1 \R_reg[2][10]  ( .D(n798), .CK(clk), .RN(rst_n), .Q(R2[10]), .QN(n542) );
  DFFRX1 \R_reg[2][9]  ( .D(n797), .CK(clk), .RN(rst_n), .Q(R2[9]), .QN(n541)
         );
  DFFRX1 \R_reg[2][6]  ( .D(n794), .CK(clk), .RN(rst_n), .Q(R2[6]), .QN(n538)
         );
  DFFRX1 \R_reg[2][5]  ( .D(n793), .CK(clk), .RN(rst_n), .Q(R2[5]), .QN(n537)
         );
  DFFRX1 \R_reg[2][0]  ( .D(n788), .CK(clk), .RN(rst_n), .Q(R2[0]), .QN(n532)
         );
  DFFRX1 \R_reg[6][15]  ( .D(n739), .CK(clk), .RN(rst_n), .Q(R6[15]), .QN(n483) );
  DFFRX1 \R_reg[6][14]  ( .D(n738), .CK(clk), .RN(rst_n), .Q(R6[14]), .QN(n482) );
  DFFRX1 \R_reg[6][13]  ( .D(n737), .CK(clk), .RN(rst_n), .Q(R6[13]), .QN(n481) );
  DFFRX1 \R_reg[6][12]  ( .D(n736), .CK(clk), .RN(rst_n), .Q(R6[12]), .QN(n480) );
  DFFRX1 \R_reg[6][11]  ( .D(n735), .CK(clk), .RN(rst_n), .Q(R6[11]), .QN(n479) );
  DFFRX1 \R_reg[6][10]  ( .D(n734), .CK(clk), .RN(rst_n), .Q(R6[10]), .QN(n478) );
  DFFRX1 \R_reg[6][9]  ( .D(n733), .CK(clk), .RN(rst_n), .Q(R6[9]), .QN(n477)
         );
  DFFRX1 \R_reg[6][8]  ( .D(n732), .CK(clk), .RN(rst_n), .Q(R6[8]), .QN(n476)
         );
  DFFRX1 \R_reg[6][7]  ( .D(n731), .CK(clk), .RN(rst_n), .Q(R6[7]), .QN(n475)
         );
  DFFRX1 \R_reg[6][6]  ( .D(n730), .CK(clk), .RN(rst_n), .Q(R6[6]), .QN(n474)
         );
  DFFRX1 \R_reg[6][5]  ( .D(n729), .CK(clk), .RN(rst_n), .Q(R6[5]), .QN(n473)
         );
  DFFRX1 \R_reg[6][0]  ( .D(n724), .CK(clk), .RN(rst_n), .Q(R6[0]), .QN(n468)
         );
  DFFRX1 \R_reg[10][15]  ( .D(n675), .CK(clk), .RN(rst_n), .Q(R10[15]), .QN(
        n419) );
  DFFRX1 \R_reg[10][14]  ( .D(n674), .CK(clk), .RN(rst_n), .Q(R10[14]), .QN(
        n418) );
  DFFRX1 \R_reg[10][13]  ( .D(n673), .CK(clk), .RN(rst_n), .Q(R10[13]), .QN(
        n417) );
  DFFRX1 \R_reg[10][12]  ( .D(n672), .CK(clk), .RN(rst_n), .Q(R10[12]), .QN(
        n416) );
  DFFRX1 \R_reg[10][11]  ( .D(n671), .CK(clk), .RN(rst_n), .Q(R10[11]), .QN(
        n415) );
  DFFRX1 \R_reg[10][10]  ( .D(n670), .CK(clk), .RN(rst_n), .Q(R10[10]), .QN(
        n414) );
  DFFRX1 \R_reg[10][9]  ( .D(n669), .CK(clk), .RN(rst_n), .Q(R10[9]), .QN(n413) );
  DFFRX1 \R_reg[10][6]  ( .D(n666), .CK(clk), .RN(rst_n), .Q(R10[6]), .QN(n410) );
  DFFRX1 \R_reg[10][5]  ( .D(n665), .CK(clk), .RN(rst_n), .Q(R10[5]), .QN(n409) );
  DFFRX1 \R_reg[10][0]  ( .D(n660), .CK(clk), .RN(rst_n), .Q(R10[0]), .QN(n404) );
  DFFRX1 \R_reg[14][15]  ( .D(n611), .CK(clk), .RN(rst_n), .Q(R14[15]), .QN(
        n355) );
  DFFRX1 \R_reg[14][14]  ( .D(n610), .CK(clk), .RN(rst_n), .Q(R14[14]), .QN(
        n354) );
  DFFRX1 \R_reg[14][13]  ( .D(n609), .CK(clk), .RN(rst_n), .Q(R14[13]), .QN(
        n353) );
  DFFRX1 \R_reg[14][12]  ( .D(n608), .CK(clk), .RN(rst_n), .Q(R14[12]), .QN(
        n352) );
  DFFRX1 \R_reg[14][11]  ( .D(n607), .CK(clk), .RN(rst_n), .Q(R14[11]), .QN(
        n351) );
  DFFRX1 \R_reg[14][10]  ( .D(n606), .CK(clk), .RN(rst_n), .Q(R14[10]), .QN(
        n350) );
  DFFRX1 \R_reg[14][9]  ( .D(n605), .CK(clk), .RN(rst_n), .Q(R14[9]), .QN(n349) );
  DFFRX1 \R_reg[14][8]  ( .D(n604), .CK(clk), .RN(rst_n), .Q(R14[8]), .QN(n348) );
  DFFRX1 \R_reg[14][7]  ( .D(n603), .CK(clk), .RN(rst_n), .Q(R14[7]), .QN(n347) );
  DFFRX1 \R_reg[14][6]  ( .D(n602), .CK(clk), .RN(rst_n), .Q(R14[6]), .QN(n346) );
  DFFRX1 \R_reg[14][5]  ( .D(n601), .CK(clk), .RN(rst_n), .Q(R14[5]), .QN(n345) );
  DFFRX1 \R_reg[14][0]  ( .D(n596), .CK(clk), .RN(rst_n), .Q(R14[0]), .QN(n340) );
  DFFRX1 \R_reg[3][8]  ( .D(n780), .CK(clk), .RN(rst_n), .Q(R3[8]), .QN(n524)
         );
  DFFRX1 \R_reg[3][7]  ( .D(n779), .CK(clk), .RN(rst_n), .Q(R3[7]), .QN(n523)
         );
  DFFRX1 \R_reg[3][4]  ( .D(n776), .CK(clk), .RN(rst_n), .Q(R3[4]), .QN(n520)
         );
  DFFRX1 \R_reg[3][3]  ( .D(n775), .CK(clk), .RN(rst_n), .Q(R3[3]), .QN(n519)
         );
  DFFRX1 \R_reg[3][2]  ( .D(n774), .CK(clk), .RN(rst_n), .Q(R3[2]), .QN(n518)
         );
  DFFRX1 \R_reg[3][1]  ( .D(n773), .CK(clk), .RN(rst_n), .Q(R3[1]), .QN(n517)
         );
  DFFRX1 \R_reg[7][4]  ( .D(n712), .CK(clk), .RN(rst_n), .Q(R7[4]), .QN(n456)
         );
  DFFRX1 \R_reg[7][3]  ( .D(n711), .CK(clk), .RN(rst_n), .Q(R7[3]), .QN(n455)
         );
  DFFRX1 \R_reg[7][2]  ( .D(n710), .CK(clk), .RN(rst_n), .Q(R7[2]), .QN(n454)
         );
  DFFRX1 \R_reg[7][1]  ( .D(n709), .CK(clk), .RN(rst_n), .Q(R7[1]), .QN(n453)
         );
  DFFRX1 \R_reg[11][8]  ( .D(n652), .CK(clk), .RN(rst_n), .Q(R11[8]), .QN(n396) );
  DFFRX1 \R_reg[11][7]  ( .D(n651), .CK(clk), .RN(rst_n), .Q(R11[7]), .QN(n395) );
  DFFRX1 \R_reg[11][4]  ( .D(n648), .CK(clk), .RN(rst_n), .Q(R11[4]), .QN(n392) );
  DFFRX1 \R_reg[11][3]  ( .D(n647), .CK(clk), .RN(rst_n), .Q(R11[3]), .QN(n391) );
  DFFRX1 \R_reg[11][2]  ( .D(n646), .CK(clk), .RN(rst_n), .Q(R11[2]), .QN(n390) );
  DFFRX1 \R_reg[11][1]  ( .D(n645), .CK(clk), .RN(rst_n), .Q(R11[1]), .QN(n389) );
  DFFRX1 \R_reg[15][4]  ( .D(n584), .CK(clk), .RN(rst_n), .Q(R15[4]), .QN(n328) );
  DFFRX1 \R_reg[15][3]  ( .D(n583), .CK(clk), .RN(rst_n), .Q(R15[3]), .QN(n327) );
  DFFRX1 \R_reg[15][2]  ( .D(n582), .CK(clk), .RN(rst_n), .Q(R15[2]), .QN(n326) );
  DFFRX1 \R_reg[15][1]  ( .D(n581), .CK(clk), .RN(rst_n), .Q(R15[1]), .QN(n325) );
  DFFRX1 \R_reg[1][8]  ( .D(n812), .CK(clk), .RN(rst_n), .Q(R1[8]), .QN(n556)
         );
  DFFRX1 \R_reg[1][7]  ( .D(n811), .CK(clk), .RN(rst_n), .Q(R1[7]), .QN(n555)
         );
  DFFRX1 \R_reg[1][4]  ( .D(n808), .CK(clk), .RN(rst_n), .Q(R1[4]), .QN(n552)
         );
  DFFRX1 \R_reg[1][3]  ( .D(n807), .CK(clk), .RN(rst_n), .Q(R1[3]), .QN(n551)
         );
  DFFRX1 \R_reg[1][2]  ( .D(n806), .CK(clk), .RN(rst_n), .Q(R1[2]), .QN(n550)
         );
  DFFRX1 \R_reg[1][1]  ( .D(n805), .CK(clk), .RN(rst_n), .Q(R1[1]), .QN(n549)
         );
  DFFRX1 \R_reg[5][8]  ( .D(n748), .CK(clk), .RN(rst_n), .Q(R5[8]), .QN(n492)
         );
  DFFRX1 \R_reg[5][7]  ( .D(n747), .CK(clk), .RN(rst_n), .Q(R5[7]), .QN(n491)
         );
  DFFRX1 \R_reg[5][4]  ( .D(n744), .CK(clk), .RN(rst_n), .Q(R5[4]), .QN(n488)
         );
  DFFRX1 \R_reg[5][3]  ( .D(n743), .CK(clk), .RN(rst_n), .Q(R5[3]), .QN(n487)
         );
  DFFRX1 \R_reg[5][2]  ( .D(n742), .CK(clk), .RN(rst_n), .Q(R5[2]), .QN(n486)
         );
  DFFRX1 \R_reg[5][1]  ( .D(n741), .CK(clk), .RN(rst_n), .Q(R5[1]), .QN(n485)
         );
  DFFRX1 \R_reg[9][8]  ( .D(n684), .CK(clk), .RN(rst_n), .Q(R9[8]), .QN(n428)
         );
  DFFRX1 \R_reg[9][7]  ( .D(n683), .CK(clk), .RN(rst_n), .Q(R9[7]), .QN(n427)
         );
  DFFRX1 \R_reg[9][4]  ( .D(n680), .CK(clk), .RN(rst_n), .Q(R9[4]), .QN(n424)
         );
  DFFRX1 \R_reg[9][3]  ( .D(n679), .CK(clk), .RN(rst_n), .Q(R9[3]), .QN(n423)
         );
  DFFRX1 \R_reg[9][2]  ( .D(n678), .CK(clk), .RN(rst_n), .Q(R9[2]), .QN(n422)
         );
  DFFRX1 \R_reg[9][1]  ( .D(n677), .CK(clk), .RN(rst_n), .Q(R9[1]), .QN(n421)
         );
  DFFRX1 \R_reg[13][8]  ( .D(n620), .CK(clk), .RN(rst_n), .Q(R13[8]), .QN(n364) );
  DFFRX1 \R_reg[13][7]  ( .D(n619), .CK(clk), .RN(rst_n), .Q(R13[7]), .QN(n363) );
  DFFRX1 \R_reg[13][4]  ( .D(n616), .CK(clk), .RN(rst_n), .Q(R13[4]), .QN(n360) );
  DFFRX1 \R_reg[13][3]  ( .D(n615), .CK(clk), .RN(rst_n), .Q(R13[3]), .QN(n359) );
  DFFRX1 \R_reg[13][2]  ( .D(n614), .CK(clk), .RN(rst_n), .Q(R13[2]), .QN(n358) );
  DFFRX1 \R_reg[13][1]  ( .D(n613), .CK(clk), .RN(rst_n), .Q(R13[1]), .QN(n357) );
  DFFRX1 \R_reg[0][8]  ( .D(n828), .CK(clk), .RN(rst_n), .Q(R0[8]), .QN(n572)
         );
  DFFRX1 \R_reg[0][7]  ( .D(n827), .CK(clk), .RN(rst_n), .Q(R0[7]), .QN(n571)
         );
  DFFRX1 \R_reg[0][4]  ( .D(n824), .CK(clk), .RN(rst_n), .Q(R0[4]), .QN(n568)
         );
  DFFRX1 \R_reg[0][3]  ( .D(n823), .CK(clk), .RN(rst_n), .Q(R0[3]), .QN(n567)
         );
  DFFRX1 \R_reg[0][2]  ( .D(n822), .CK(clk), .RN(rst_n), .Q(R0[2]), .QN(n566)
         );
  DFFRX1 \R_reg[0][1]  ( .D(n821), .CK(clk), .RN(rst_n), .Q(R0[1]), .QN(n565)
         );
  DFFRX1 \R_reg[4][8]  ( .D(n764), .CK(clk), .RN(rst_n), .Q(R4[8]), .QN(n508)
         );
  DFFRX1 \R_reg[4][7]  ( .D(n763), .CK(clk), .RN(rst_n), .Q(R4[7]), .QN(n507)
         );
  DFFRX1 \R_reg[4][4]  ( .D(n760), .CK(clk), .RN(rst_n), .Q(R4[4]), .QN(n504)
         );
  DFFRX1 \R_reg[4][3]  ( .D(n759), .CK(clk), .RN(rst_n), .Q(R4[3]), .QN(n503)
         );
  DFFRX1 \R_reg[4][2]  ( .D(n758), .CK(clk), .RN(rst_n), .Q(R4[2]), .QN(n502)
         );
  DFFRX1 \R_reg[4][1]  ( .D(n757), .CK(clk), .RN(rst_n), .Q(R4[1]), .QN(n501)
         );
  DFFRX1 \R_reg[8][8]  ( .D(n700), .CK(clk), .RN(rst_n), .Q(R8[8]), .QN(n444)
         );
  DFFRX1 \R_reg[8][7]  ( .D(n699), .CK(clk), .RN(rst_n), .Q(R8[7]), .QN(n443)
         );
  DFFRX1 \R_reg[8][4]  ( .D(n696), .CK(clk), .RN(rst_n), .Q(R8[4]), .QN(n440)
         );
  DFFRX1 \R_reg[8][3]  ( .D(n695), .CK(clk), .RN(rst_n), .Q(R8[3]), .QN(n439)
         );
  DFFRX1 \R_reg[8][2]  ( .D(n694), .CK(clk), .RN(rst_n), .Q(R8[2]), .QN(n438)
         );
  DFFRX1 \R_reg[8][1]  ( .D(n693), .CK(clk), .RN(rst_n), .Q(R8[1]), .QN(n437)
         );
  DFFRX1 \R_reg[12][8]  ( .D(n636), .CK(clk), .RN(rst_n), .Q(R12[8]), .QN(n380) );
  DFFRX1 \R_reg[12][7]  ( .D(n635), .CK(clk), .RN(rst_n), .Q(R12[7]), .QN(n379) );
  DFFRX1 \R_reg[12][4]  ( .D(n632), .CK(clk), .RN(rst_n), .Q(R12[4]), .QN(n376) );
  DFFRX1 \R_reg[12][3]  ( .D(n631), .CK(clk), .RN(rst_n), .Q(R12[3]), .QN(n375) );
  DFFRX1 \R_reg[12][2]  ( .D(n630), .CK(clk), .RN(rst_n), .Q(R12[2]), .QN(n374) );
  DFFRX1 \R_reg[12][1]  ( .D(n629), .CK(clk), .RN(rst_n), .Q(R12[1]), .QN(n373) );
  DFFRX1 \R_reg[2][8]  ( .D(n796), .CK(clk), .RN(rst_n), .Q(R2[8]), .QN(n540)
         );
  DFFRX1 \R_reg[2][7]  ( .D(n795), .CK(clk), .RN(rst_n), .Q(R2[7]), .QN(n539)
         );
  DFFRX1 \R_reg[2][4]  ( .D(n792), .CK(clk), .RN(rst_n), .Q(R2[4]), .QN(n536)
         );
  DFFRX1 \R_reg[2][3]  ( .D(n791), .CK(clk), .RN(rst_n), .Q(R2[3]), .QN(n535)
         );
  DFFRX1 \R_reg[2][2]  ( .D(n790), .CK(clk), .RN(rst_n), .Q(R2[2]), .QN(n534)
         );
  DFFRX1 \R_reg[2][1]  ( .D(n789), .CK(clk), .RN(rst_n), .Q(R2[1]), .QN(n533)
         );
  DFFRX1 \R_reg[6][4]  ( .D(n728), .CK(clk), .RN(rst_n), .Q(R6[4]), .QN(n472)
         );
  DFFRX1 \R_reg[6][3]  ( .D(n727), .CK(clk), .RN(rst_n), .Q(R6[3]), .QN(n471)
         );
  DFFRX1 \R_reg[6][2]  ( .D(n726), .CK(clk), .RN(rst_n), .Q(R6[2]), .QN(n470)
         );
  DFFRX1 \R_reg[6][1]  ( .D(n725), .CK(clk), .RN(rst_n), .Q(R6[1]), .QN(n469)
         );
  DFFRX1 \R_reg[10][8]  ( .D(n668), .CK(clk), .RN(rst_n), .Q(R10[8]), .QN(n412) );
  DFFRX1 \R_reg[10][7]  ( .D(n667), .CK(clk), .RN(rst_n), .Q(R10[7]), .QN(n411) );
  DFFRX1 \R_reg[10][4]  ( .D(n664), .CK(clk), .RN(rst_n), .Q(R10[4]), .QN(n408) );
  DFFRX1 \R_reg[10][3]  ( .D(n663), .CK(clk), .RN(rst_n), .Q(R10[3]), .QN(n407) );
  DFFRX1 \R_reg[10][2]  ( .D(n662), .CK(clk), .RN(rst_n), .Q(R10[2]), .QN(n406) );
  DFFRX1 \R_reg[10][1]  ( .D(n661), .CK(clk), .RN(rst_n), .Q(R10[1]), .QN(n405) );
  DFFRX1 \R_reg[14][4]  ( .D(n600), .CK(clk), .RN(rst_n), .Q(R14[4]), .QN(n344) );
  DFFRX1 \R_reg[14][3]  ( .D(n599), .CK(clk), .RN(rst_n), .Q(R14[3]), .QN(n343) );
  DFFRX1 \R_reg[14][2]  ( .D(n598), .CK(clk), .RN(rst_n), .Q(R14[2]), .QN(n342) );
  DFFRX1 \R_reg[14][1]  ( .D(n597), .CK(clk), .RN(rst_n), .Q(R14[1]), .QN(n341) );
  CLKINVX3 U609 ( .A(n1349), .Y(MUXB[13]) );
  NAND2XL U610 ( .A(n1421), .B(n1520), .Y(n1214) );
  NAND2XL U611 ( .A(n1423), .B(n1520), .Y(n1283) );
  NAND2XL U612 ( .A(n1419), .B(n1520), .Y(n1252) );
  NOR2XL U613 ( .A(n1520), .B(n874), .Y(n1524) );
  CLKINVX1 U614 ( .A(n1475), .Y(n1448) );
  NOR2XL U615 ( .A(n1323), .B(n857), .Y(n1274) );
  MXI2XL U616 ( .A(n1323), .B(n1406), .S0(N201), .Y(n1234) );
  NOR2XL U617 ( .A(n1323), .B(n874), .Y(n1324) );
  NAND2XL U618 ( .A(N201), .B(n1323), .Y(n1277) );
  MXI2X2 U619 ( .A(N101), .B(constant[14]), .S0(control[13]), .Y(n1323) );
  MXI2X1 U620 ( .A(N114), .B(constant[1]), .S0(control[13]), .Y(n1515) );
  MXI4X1 U621 ( .A(n1005), .B(n1006), .C(n1007), .D(n1008), .S0(N60), .S1(N59), 
        .Y(N114) );
  MXI2X2 U622 ( .A(N113), .B(constant[2]), .S0(control[13]), .Y(n1522) );
  MXI4X1 U623 ( .A(n1009), .B(n1010), .C(n1011), .D(n1012), .S0(N60), .S1(N59), 
        .Y(N113) );
  MXI2X2 U624 ( .A(N112), .B(constant[3]), .S0(control[13]), .Y(n1521) );
  MXI4X2 U625 ( .A(n1013), .B(n1014), .C(n1015), .D(n1016), .S0(N60), .S1(N59), 
        .Y(N112) );
  MXI4X1 U626 ( .A(R8[3]), .B(R9[3]), .C(R10[3]), .D(R11[3]), .S0(N57), .S1(
        n1066), .Y(n1014) );
  MXI4X1 U627 ( .A(R0[3]), .B(R1[3]), .C(R2[3]), .D(R3[3]), .S0(N57), .S1(
        n1066), .Y(n1013) );
  MXI2X2 U628 ( .A(N111), .B(constant[4]), .S0(control[13]), .Y(n1520) );
  MXI4X1 U629 ( .A(n1017), .B(n1018), .C(n1019), .D(n1020), .S0(N60), .S1(N59), 
        .Y(N111) );
  MXI4X1 U630 ( .A(R8[4]), .B(R9[4]), .C(R10[4]), .D(R11[4]), .S0(N57), .S1(
        n1067), .Y(n1018) );
  MXI4X1 U631 ( .A(R0[4]), .B(R1[4]), .C(R2[4]), .D(R3[4]), .S0(N57), .S1(
        n1067), .Y(n1017) );
  MXI2X2 U632 ( .A(N110), .B(constant[5]), .S0(control[13]), .Y(n1474) );
  AND2X2 U633 ( .A(n1856), .B(n1602), .Y(n876) );
  AND2X2 U634 ( .A(n1856), .B(n1584), .Y(n877) );
  AND2X2 U635 ( .A(n1856), .B(n1657), .Y(n878) );
  AND2X2 U636 ( .A(n1856), .B(n1640), .Y(n879) );
  CLKINVX1 U637 ( .A(control[3]), .Y(n1287) );
  MXI2X2 U638 ( .A(n868), .B(constant[7]), .S0(control[13]), .Y(n1422) );
  MXI4X1 U639 ( .A(n1029), .B(n1030), .C(n1031), .D(n1032), .S0(N60), .S1(N59), 
        .Y(n868) );
  MXI4X1 U640 ( .A(R12[7]), .B(R13[7]), .C(R14[7]), .D(R15[7]), .S0(N57), .S1(
        n1068), .Y(n1032) );
  MXI4X1 U641 ( .A(R4[7]), .B(R5[7]), .C(R6[7]), .D(R7[7]), .S0(N57), .S1(
        n1068), .Y(n1031) );
  MXI2X1 U642 ( .A(N103), .B(constant[12]), .S0(control[13]), .Y(n1346) );
  NAND2X1 U643 ( .A(N201), .B(n1287), .Y(n857) );
  NAND2X1 U644 ( .A(n1328), .B(n1179), .Y(N203) );
  MXI2X1 U645 ( .A(N102), .B(constant[13]), .S0(control[13]), .Y(n1349) );
  MXI4X1 U646 ( .A(n1053), .B(n1054), .C(n1055), .D(n1056), .S0(N60), .S1(N59), 
        .Y(N102) );
  MX4X1 U647 ( .A(n1061), .B(n1062), .C(n1063), .D(n1064), .S0(N60), .S1(N59), 
        .Y(n872) );
  AND2X2 U648 ( .A(N504), .B(n901), .Y(n1783) );
  MXI2X2 U649 ( .A(N107), .B(constant[8]), .S0(control[13]), .Y(n1418) );
  MXI4X1 U650 ( .A(n1033), .B(n1034), .C(n1035), .D(n1036), .S0(N60), .S1(N59), 
        .Y(N107) );
  MXI2X2 U651 ( .A(N106), .B(constant[9]), .S0(control[13]), .Y(n1420) );
  MXI2X1 U652 ( .A(N105), .B(constant[10]), .S0(control[13]), .Y(n1347) );
  NAND2X1 U653 ( .A(n840), .B(n1536), .Y(BUSB[1]) );
  NAND4X1 U654 ( .A(n1512), .B(n1511), .C(n1510), .D(n1509), .Y(BUSB[2]) );
  AO21X1 U655 ( .A0(n1489), .A1(n1488), .B0(n1487), .Y(n855) );
  NAND4X1 U656 ( .A(n1470), .B(n1469), .C(n1468), .D(n1467), .Y(BUSB[4]) );
  NAND4X1 U657 ( .A(n1454), .B(n1453), .C(n1452), .D(n1451), .Y(BUSB[5]) );
  NAND4BBXL U658 ( .AN(n853), .BN(n854), .C(n1433), .D(n1432), .Y(BUSB[6]) );
  MXI4X1 U659 ( .A(n1077), .B(n1078), .C(n1079), .D(n1080), .S0(N64), .S1(N63), 
        .Y(BUSA[1]) );
  MXI4X1 U660 ( .A(n1081), .B(n1082), .C(n1083), .D(n1084), .S0(N64), .S1(N63), 
        .Y(BUSA[2]) );
  MXI4X1 U661 ( .A(n1085), .B(n1086), .C(n1087), .D(n1088), .S0(N64), .S1(N63), 
        .Y(BUSA[3]) );
  MXI4X1 U662 ( .A(n1089), .B(n1090), .C(n1091), .D(n1092), .S0(N64), .S1(N63), 
        .Y(BUSA[4]) );
  MXI4X1 U663 ( .A(n1093), .B(n1094), .C(n1095), .D(n1096), .S0(N64), .S1(N63), 
        .Y(BUSA[5]) );
  MXI4X1 U664 ( .A(n1097), .B(n1098), .C(n1099), .D(n1100), .S0(N64), .S1(N63), 
        .Y(BUSA[6]) );
  MXI4X1 U665 ( .A(n1101), .B(n1102), .C(n1103), .D(n1104), .S0(N64), .S1(N63), 
        .Y(BUSA[7]) );
  OA21XL U666 ( .A0(n1862), .A1(n1834), .B0(n1833), .Y(n837) );
  OA21XL U667 ( .A0(n1717), .A1(n1834), .B0(n1716), .Y(n838) );
  OR2X1 U668 ( .A(n1838), .B(n1837), .Y(n839) );
  AND3X2 U669 ( .A(n1534), .B(n1537), .C(n1535), .Y(n840) );
  CLKINVX1 U670 ( .A(n870), .Y(n1406) );
  MXI2X1 U671 ( .A(n872), .B(n871), .S0(control[13]), .Y(n870) );
  OR2X1 U672 ( .A(n1418), .B(n869), .Y(n841) );
  OR2X1 U673 ( .A(n1347), .B(n869), .Y(n842) );
  OR2X1 U674 ( .A(n1420), .B(n869), .Y(n843) );
  AND2X2 U675 ( .A(BUSA[10]), .B(n1173), .Y(n844) );
  AND2X2 U676 ( .A(BUSA[12]), .B(n1173), .Y(n845) );
  AND2X2 U677 ( .A(BUSA[8]), .B(n1173), .Y(n846) );
  NAND3X1 U678 ( .A(n920), .B(control[12]), .C(n1551), .Y(n847) );
  CLKINVX1 U679 ( .A(n1522), .Y(MUXB[2]) );
  MXI4X1 U680 ( .A(n1021), .B(n1022), .C(n1023), .D(n1024), .S0(N60), .S1(N59), 
        .Y(N110) );
  MXI4X1 U681 ( .A(n1057), .B(n1058), .C(n1059), .D(n1060), .S0(N60), .S1(N59), 
        .Y(N101) );
  MXI4X1 U682 ( .A(n1037), .B(n1038), .C(n1039), .D(n1040), .S0(N60), .S1(N59), 
        .Y(N106) );
  INVX1 U683 ( .A(n1515), .Y(MUXB[1]) );
  XNOR2XL U684 ( .A(\FUResult[15] ), .B(BUSA[15]), .Y(n1863) );
  CLKINVX1 U685 ( .A(n1441), .Y(MUXB[6]) );
  CLKINVX1 U686 ( .A(n851), .Y(n1384) );
  MXI4X1 U687 ( .A(n1001), .B(n1002), .C(n1003), .D(n1004), .S0(N60), .S1(N59), 
        .Y(N115) );
  NAND2X1 U688 ( .A(N115), .B(n848), .Y(n849) );
  NAND2X1 U689 ( .A(n849), .B(n850), .Y(n851) );
  CLKINVX1 U690 ( .A(BUSB[0]), .Y(n1552) );
  NAND3XL U691 ( .A(n1829), .B(n1828), .C(n1827), .Y(\FUResult[15] ) );
  MXI4X1 U692 ( .A(R0[14]), .B(R1[14]), .C(R2[14]), .D(R3[14]), .S0(N57), .S1(
        n1070), .Y(n1057) );
  MXI4X1 U693 ( .A(R0[12]), .B(R1[12]), .C(R2[12]), .D(R3[12]), .S0(N57), .S1(
        n1069), .Y(n1049) );
  CLKMX2X2 U694 ( .A(N104), .B(constant[11]), .S0(control[13]), .Y(n852) );
  MXI4X1 U695 ( .A(n1045), .B(n1046), .C(n1047), .D(n1048), .S0(N60), .S1(N59), 
        .Y(N104) );
  CLKINVX1 U696 ( .A(N201), .Y(n1175) );
  NAND2X1 U697 ( .A(constant[0]), .B(control[13]), .Y(n850) );
  INVX1 U698 ( .A(control[13]), .Y(n848) );
  NAND2XL U699 ( .A(n1421), .B(n1384), .Y(n1210) );
  NAND2XL U700 ( .A(control[3]), .B(n1384), .Y(n1248) );
  MXI2XL U701 ( .A(n1515), .B(n1384), .S0(N201), .Y(n1288) );
  AND2X2 U702 ( .A(N505), .B(n901), .Y(n1804) );
  AND2X2 U703 ( .A(N466), .B(n1857), .Y(n1790) );
  INVXL U704 ( .A(BUSB[4]), .Y(n1621) );
  OA21XL U705 ( .A0(n1281), .A1(n1484), .B0(n1280), .Y(n856) );
  MXI4XL U706 ( .A(R4[9]), .B(R5[9]), .C(R6[9]), .D(R7[9]), .S0(N57), .S1(
        n1068), .Y(n1039) );
  MXI4XL U707 ( .A(R12[9]), .B(R13[9]), .C(R14[9]), .D(R15[9]), .S0(N57), .S1(
        n1068), .Y(n1040) );
  MXI4XL U708 ( .A(R4[2]), .B(R5[2]), .C(R6[2]), .D(R7[2]), .S0(N57), .S1(
        n1066), .Y(n1011) );
  MXI4XL U709 ( .A(R12[2]), .B(R13[2]), .C(R14[2]), .D(R15[2]), .S0(N57), .S1(
        n1066), .Y(n1012) );
  MXI4XL U710 ( .A(R4[1]), .B(R5[1]), .C(R6[1]), .D(R7[1]), .S0(N57), .S1(
        n1066), .Y(n1007) );
  MXI4XL U711 ( .A(R12[1]), .B(R13[1]), .C(R14[1]), .D(R15[1]), .S0(N57), .S1(
        n1066), .Y(n1008) );
  MXI4XL U712 ( .A(R0[1]), .B(R1[1]), .C(R2[1]), .D(R3[1]), .S0(N57), .S1(
        n1066), .Y(n1005) );
  MXI4XL U713 ( .A(R8[1]), .B(R9[1]), .C(R10[1]), .D(R11[1]), .S0(N57), .S1(
        n1066), .Y(n1006) );
  MXI4XL U714 ( .A(R4[14]), .B(R5[14]), .C(R6[14]), .D(R7[14]), .S0(N57), .S1(
        n1070), .Y(n1059) );
  MXI4XL U715 ( .A(R12[14]), .B(R13[14]), .C(R14[14]), .D(R15[14]), .S0(N57), 
        .S1(n1070), .Y(n1060) );
  MXI4XL U716 ( .A(R8[13]), .B(R9[13]), .C(R10[13]), .D(R11[13]), .S0(N57), 
        .S1(n1070), .Y(n1054) );
  MXI4XL U717 ( .A(R8[6]), .B(R9[6]), .C(R10[6]), .D(R11[6]), .S0(N57), .S1(
        n1067), .Y(n1026) );
  MXI4XL U718 ( .A(R8[14]), .B(R9[14]), .C(R10[14]), .D(R11[14]), .S0(N57), 
        .S1(n1070), .Y(n1058) );
  MXI4XL U719 ( .A(R0[13]), .B(R1[13]), .C(R2[13]), .D(R3[13]), .S0(N57), .S1(
        n1070), .Y(n1053) );
  MXI4XL U720 ( .A(R0[6]), .B(R1[6]), .C(R2[6]), .D(R3[6]), .S0(N57), .S1(
        n1067), .Y(n1025) );
  CLKINVX1 U721 ( .A(BUSB[8]), .Y(n1689) );
  CLKINVX1 U722 ( .A(n1162), .Y(n1348) );
  AOI21X1 U723 ( .A0(N302), .A1(n1514), .B0(n1382), .Y(n1393) );
  AOI22X1 U724 ( .A0(N299), .A1(n1514), .B0(n1450), .B1(n1498), .Y(n1451) );
  NOR3XL U725 ( .A(n1533), .B(n1532), .C(n1531), .Y(n1534) );
  NAND2XL U726 ( .A(N208), .B(n1513), .Y(n1537) );
  AOI21X1 U727 ( .A0(n1334), .A1(n1330), .B0(n1329), .Y(n1483) );
  NOR2XL U728 ( .A(n1384), .B(n1405), .Y(n1385) );
  NAND2X1 U729 ( .A(n1457), .B(n1388), .Y(n1199) );
  NAND2XL U730 ( .A(n1421), .B(n1349), .Y(n1352) );
  NOR4X1 U731 ( .A(n1826), .B(n897), .C(n1825), .D(n1824), .Y(n1827) );
  NAND2BX1 U732 ( .AN(n1482), .B(n1484), .Y(n1456) );
  NOR2X1 U733 ( .A(n1322), .B(n1321), .Y(n1327) );
  NAND2X1 U734 ( .A(n1203), .B(n1184), .Y(n1482) );
  NAND2X1 U735 ( .A(n1175), .B(n1287), .Y(n1444) );
  CLKINVX1 U736 ( .A(n1347), .Y(MUXB[10]) );
  MXI4X1 U737 ( .A(R12[5]), .B(R13[5]), .C(R14[5]), .D(R15[5]), .S0(N57), .S1(
        n1067), .Y(n1024) );
  MXI4X1 U738 ( .A(R4[5]), .B(R5[5]), .C(R6[5]), .D(R7[5]), .S0(N57), .S1(
        n1067), .Y(n1023) );
  MXI4X1 U739 ( .A(R0[2]), .B(R1[2]), .C(R2[2]), .D(R3[2]), .S0(N57), .S1(
        n1066), .Y(n1009) );
  MXI4X1 U740 ( .A(R0[8]), .B(R1[8]), .C(R2[8]), .D(R3[8]), .S0(N57), .S1(
        n1068), .Y(n1033) );
  MXI4X1 U741 ( .A(R0[9]), .B(R1[9]), .C(R2[9]), .D(R3[9]), .S0(N57), .S1(
        n1068), .Y(n1037) );
  MXI4X1 U742 ( .A(R0[5]), .B(R1[5]), .C(R2[5]), .D(R3[5]), .S0(N57), .S1(
        n1067), .Y(n1021) );
  MXI4X1 U743 ( .A(R8[2]), .B(R9[2]), .C(R10[2]), .D(R11[2]), .S0(N57), .S1(
        n1066), .Y(n1010) );
  MXI4X1 U744 ( .A(R8[8]), .B(R9[8]), .C(R10[8]), .D(R11[8]), .S0(N57), .S1(
        n1068), .Y(n1034) );
  MXI4X1 U745 ( .A(R8[9]), .B(R9[9]), .C(R10[9]), .D(R11[9]), .S0(N57), .S1(
        n1068), .Y(n1038) );
  MXI4X1 U746 ( .A(R8[5]), .B(R9[5]), .C(R10[5]), .D(R11[5]), .S0(N57), .S1(
        n1067), .Y(n1022) );
  MXI4X1 U747 ( .A(R8[12]), .B(R9[12]), .C(R10[12]), .D(R11[12]), .S0(N57), 
        .S1(n1069), .Y(n1050) );
  CLKINVX1 U748 ( .A(constant[15]), .Y(n871) );
  BUFX4 U749 ( .A(N58), .Y(n1072) );
  CLKINVX1 U750 ( .A(control[4]), .Y(n1330) );
  BUFX2 U751 ( .A(N58), .Y(n1071) );
  NOR2XL U752 ( .A(n1347), .B(n873), .Y(n1300) );
  NOR2XL U753 ( .A(n1347), .B(n857), .Y(n1367) );
  NOR2XL U754 ( .A(n1347), .B(n874), .Y(n1400) );
  NOR2XL U755 ( .A(n1347), .B(n1163), .Y(n1256) );
  INVXL U756 ( .A(BUSB[7]), .Y(n1673) );
  INVXL U757 ( .A(BUSB[9]), .Y(n1707) );
  NOR2XL U758 ( .A(n1529), .B(n1475), .Y(n1377) );
  NOR2XL U759 ( .A(n1459), .B(n1475), .Y(n1389) );
  NOR2BXL U760 ( .AN(n1434), .B(n1526), .Y(n1437) );
  NOR2XL U761 ( .A(n1459), .B(n1526), .Y(n1460) );
  NOR2XL U762 ( .A(n1458), .B(n1528), .Y(n1461) );
  INVX1 U763 ( .A(n1388), .Y(n1459) );
  INVX1 U764 ( .A(n1434), .Y(n1529) );
  NAND2XL U765 ( .A(n1759), .B(BUSB[7]), .Y(n1671) );
  OR3X2 U766 ( .A(n1417), .B(n1416), .C(n1490), .Y(n853) );
  AO21XL U767 ( .A0(n1457), .A1(n1500), .B0(n1428), .Y(n854) );
  NOR3XL U768 ( .A(n1391), .B(n1390), .C(n1389), .Y(n1392) );
  NOR3XL U769 ( .A(n1438), .B(n1437), .C(n1436), .Y(n1454) );
  AOI21XL U770 ( .A0(N212), .A1(n1513), .B0(n1449), .Y(n1452) );
  NAND2XL U771 ( .A(n1498), .B(n1396), .Y(n1413) );
  NOR2XL U772 ( .A(n1410), .B(n1409), .Y(n1411) );
  AOI21XL U773 ( .A0(N214), .A1(n1513), .B0(n1397), .Y(n1412) );
  AOI21XL U774 ( .A0(N303), .A1(n1514), .B0(n1363), .Y(n1379) );
  NOR2XL U775 ( .A(n1491), .B(n1517), .Y(n1492) );
  NAND2X1 U776 ( .A(N296), .B(n1514), .Y(n1511) );
  AOI21X1 U777 ( .A0(N300), .A1(n1514), .B0(n1431), .Y(n1432) );
  NAND2XL U778 ( .A(N216), .B(n1513), .Y(n1380) );
  NAND2X1 U779 ( .A(N295), .B(n1514), .Y(n1536) );
  NOR2XL U780 ( .A(n1435), .B(n1371), .Y(n1375) );
  NOR2XL U781 ( .A(n1258), .B(n1241), .Y(n1197) );
  NOR2XL U782 ( .A(n1305), .B(n1300), .Y(n1198) );
  NOR2XL U783 ( .A(n1526), .B(n1505), .Y(n1417) );
  NOR2XL U784 ( .A(n1504), .B(n1475), .Y(n1428) );
  NOR2XL U785 ( .A(n1435), .B(n1430), .Y(n1357) );
  NOR2XL U786 ( .A(n1387), .B(n1435), .Y(n1390) );
  INVXL U787 ( .A(n1471), .Y(n1865) );
  NAND2BX1 U788 ( .AN(n1735), .B(n1723), .Y(n1724) );
  NOR2XL U789 ( .A(n1517), .B(n1516), .Y(n1518) );
  NAND2XL U790 ( .A(N301), .B(n1514), .Y(n1414) );
  NOR2XL U791 ( .A(n1367), .B(n1366), .Y(n1368) );
  NOR2XL U792 ( .A(n1365), .B(n1364), .Y(n1369) );
  NAND2XL U793 ( .A(N215), .B(n1513), .Y(n1394) );
  INVX1 U794 ( .A(n1334), .Y(n1486) );
  NAND2BXL U795 ( .AN(n1435), .B(n1381), .Y(n1314) );
  NAND2BXL U796 ( .AN(n1526), .B(n1478), .Y(n1479) );
  INVX1 U797 ( .A(n1316), .Y(n1458) );
  INVX1 U798 ( .A(N467), .Y(n1810) );
  NAND2BX1 U799 ( .AN(n1773), .B(n1761), .Y(n1762) );
  INVXL U800 ( .A(n1442), .Y(n1443) );
  NOR3XL U801 ( .A(n1400), .B(n1325), .C(n1364), .Y(n1282) );
  MXI2XL U802 ( .A(n1760), .B(n1759), .S0(n1552), .Y(n1553) );
  NAND2XL U803 ( .A(n1800), .B(BUSB[0]), .Y(n1563) );
  NOR3XL U804 ( .A(n1366), .B(n1321), .C(n1274), .Y(n1226) );
  NAND2XL U805 ( .A(n1759), .B(BUSB[4]), .Y(n1619) );
  NAND2XL U806 ( .A(n1498), .B(n1244), .Y(n1245) );
  NAND2XL U807 ( .A(n1238), .B(n1500), .Y(n1246) );
  NAND2BX1 U808 ( .AN(n1701), .B(n1690), .Y(n1691) );
  INVXL U809 ( .A(n1241), .Y(n1242) );
  CLKINVX1 U810 ( .A(n1823), .Y(n1759) );
  NAND4BBXL U811 ( .AN(n1320), .BN(n1336), .C(n1319), .D(n1318), .Y(BUSB[12])
         );
  AOI21XL U812 ( .A0(n1385), .A1(n1464), .B0(n1415), .Y(n1386) );
  AOI21XL U813 ( .A0(n1407), .A1(n1482), .B0(n1415), .Y(n1408) );
  NAND2XL U814 ( .A(n1419), .B(n1515), .Y(n1212) );
  NAND2XL U815 ( .A(n1348), .B(n1521), .Y(n1211) );
  CLKINVX1 U816 ( .A(n1223), .Y(n1514) );
  INVXL U817 ( .A(n1300), .Y(n1301) );
  NAND2XL U818 ( .A(n1423), .B(n1441), .Y(n1213) );
  NAND2XL U819 ( .A(n1348), .B(n1422), .Y(n1215) );
  NAND2XL U820 ( .A(n1348), .B(n1347), .Y(n1353) );
  NAND4BBX2 U821 ( .AN(n1495), .BN(n855), .C(n1494), .D(n1493), .Y(BUSB[3]) );
  INVX1 U822 ( .A(n1203), .Y(n1513) );
  NOR3XL U823 ( .A(n1486), .B(n1335), .C(n1484), .Y(n1337) );
  NOR2XL U824 ( .A(n1349), .B(n857), .Y(n1240) );
  NAND2XL U825 ( .A(n1421), .B(n1522), .Y(n1284) );
  NAND2XL U826 ( .A(n1348), .B(n1474), .Y(n1285) );
  NAND2XL U827 ( .A(n1419), .B(n1522), .Y(n1312) );
  NAND2XL U828 ( .A(n1421), .B(n1515), .Y(n1310) );
  NAND3XL U829 ( .A(n1234), .B(n1287), .C(n1482), .Y(n1237) );
  MXI2XL U830 ( .A(n1406), .B(n1323), .S0(n1348), .Y(n1235) );
  NOR2XL U831 ( .A(n1349), .B(n873), .Y(n1321) );
  AOI2BB2XL U832 ( .B0(N515), .B1(n1852), .A0N(n1584), .A1N(n847), .Y(n1594)
         );
  NOR3XL U833 ( .A(n1182), .B(n1181), .C(n1180), .Y(n1187) );
  NOR2XL U834 ( .A(n1515), .B(n857), .Y(n1182) );
  NOR2XL U835 ( .A(n1350), .B(n1162), .Y(n1322) );
  NOR2XL U836 ( .A(n1441), .B(n874), .Y(n1472) );
  NOR2XL U837 ( .A(n1418), .B(n1162), .Y(n1305) );
  NAND2XL U838 ( .A(n869), .B(n1471), .Y(n1317) );
  AOI2BB2XL U839 ( .B0(N520), .B1(n1852), .A0N(n1673), .A1N(n847), .Y(n1683)
         );
  AOI2BB2XL U840 ( .B0(N519), .B1(n1852), .A0N(n1657), .A1N(n847), .Y(n1667)
         );
  NAND2XL U841 ( .A(n1348), .B(n1441), .Y(n1426) );
  NAND2X1 U842 ( .A(n1383), .B(n1464), .Y(n1435) );
  NOR2XL U843 ( .A(n1446), .B(n1445), .Y(n1527) );
  INVXL U844 ( .A(n1439), .Y(n1440) );
  NOR2XL U845 ( .A(n1325), .B(n1324), .Y(n1326) );
  NOR2XL U846 ( .A(n1399), .B(n1398), .Y(n1403) );
  NOR2XL U847 ( .A(n1401), .B(n1400), .Y(n1402) );
  NAND2X1 U848 ( .A(n1238), .B(n1464), .Y(n1517) );
  NAND3BX1 U849 ( .AN(n1755), .B(n1795), .C(n1756), .Y(n1763) );
  NAND2XL U850 ( .A(n1348), .B(n1349), .Y(n1278) );
  NAND2XL U851 ( .A(n1348), .B(n1520), .Y(n1311) );
  NOR2XL U852 ( .A(n1435), .B(n1496), .Y(n1416) );
  NOR2XL U853 ( .A(n1258), .B(n1257), .Y(n1259) );
  NOR2BXL U854 ( .AN(n1500), .B(n1362), .Y(n1344) );
  NOR2XL U855 ( .A(n1349), .B(n1163), .Y(n1273) );
  NOR2XL U856 ( .A(n856), .B(n1485), .Y(n1438) );
  NOR2XL U857 ( .A(n856), .B(n1362), .Y(n1363) );
  OAI2BB1XL U858 ( .A0N(n1178), .A1N(n1463), .B0(n1405), .Y(N204) );
  NOR2XL U859 ( .A(n1515), .B(n898), .Y(n1519) );
  NOR2XL U860 ( .A(n1522), .B(n898), .Y(n1497) );
  NOR2XL U861 ( .A(n1304), .B(n1188), .Y(n1191) );
  NOR2XL U862 ( .A(n1189), .B(n1257), .Y(n1190) );
  NOR2XL U863 ( .A(n1520), .B(n1162), .Y(n1188) );
  NOR2XL U864 ( .A(n1193), .B(n1192), .Y(n1196) );
  NOR2XL U865 ( .A(n1240), .B(n1194), .Y(n1195) );
  NOR2XL U866 ( .A(n1346), .B(n1162), .Y(n1193) );
  NOR2XL U867 ( .A(n1305), .B(n1304), .Y(n1308) );
  NOR2XL U868 ( .A(n1306), .B(n1502), .Y(n1307) );
  NOR2XL U869 ( .A(n1483), .B(n1331), .Y(n1332) );
  NAND2XL U870 ( .A(n1482), .B(n1463), .Y(n1331) );
  CLKINVX1 U871 ( .A(n1362), .Y(n1383) );
  NAND2XL U872 ( .A(n1423), .B(n1522), .Y(n1209) );
  OR2XL U873 ( .A(n1415), .B(n1266), .Y(n1336) );
  INVX1 U874 ( .A(n1455), .Y(n1490) );
  OR2X1 U875 ( .A(BUSA[7]), .B(\add_233/carry[7] ), .Y(\add_233/carry[8] ) );
  OR2X1 U876 ( .A(BUSA[1]), .B(BUSA[0]), .Y(\add_233/carry[2] ) );
  OR2X1 U877 ( .A(BUSA[4]), .B(\add_233/carry[4] ), .Y(\add_233/carry[5] ) );
  AND2XL U878 ( .A(n869), .B(n1471), .Y(n898) );
  NAND2X1 U879 ( .A(n1798), .B(n1797), .Y(n1847) );
  OR3X2 U880 ( .A(n1780), .B(BUSA[12]), .C(BUSA[13]), .Y(n1791) );
  AOI21XL U881 ( .A0(n1759), .A1(BUSB[8]), .B0(n1813), .Y(n1687) );
  NOR2XL U882 ( .A(n1240), .B(n1239), .Y(n1243) );
  AOI21XL U883 ( .A0(n1450), .A1(n1457), .B0(n1289), .Y(n1294) );
  NOR2XL U884 ( .A(n1530), .B(n1516), .Y(n1289) );
  NOR2XL U885 ( .A(n1491), .B(n1530), .Y(n1218) );
  NOR2XL U886 ( .A(n1602), .B(n847), .Y(n1595) );
  NOR2XL U887 ( .A(n1621), .B(n847), .Y(n1614) );
  NOR2XL U888 ( .A(n1640), .B(n847), .Y(n1633) );
  NOR2XL U889 ( .A(n1349), .B(n898), .Y(n1272) );
  NOR2XL U890 ( .A(n1264), .B(n1317), .Y(n1208) );
  NOR2XL U891 ( .A(n1485), .B(n1430), .Y(n1253) );
  NOR2XL U892 ( .A(n1323), .B(n898), .Y(n1233) );
  NOR2XL U893 ( .A(n1530), .B(n1496), .Y(n1254) );
  MXI2XL U894 ( .A(n1760), .B(n1759), .S0(n1602), .Y(n1603) );
  MXI2XL U895 ( .A(n1760), .B(n1759), .S0(n1621), .Y(n1622) );
  MXI2XL U896 ( .A(n1760), .B(n1759), .S0(n1673), .Y(n1674) );
  MXI2XL U897 ( .A(n1760), .B(n1759), .S0(n1640), .Y(n1641) );
  MXI2XL U898 ( .A(n1760), .B(n1759), .S0(n1584), .Y(n1585) );
  MXI2XL U899 ( .A(n1760), .B(n1759), .S0(n1657), .Y(n1658) );
  AOI21XL U900 ( .A0(n128), .A1(n1840), .B0(n859), .Y(n858) );
  AO21X1 U901 ( .A0(N68), .A1(n1868), .B0(n1809), .Y(n859) );
  CLKINVX1 U902 ( .A(n1539), .Y(n1852) );
  NAND2X1 U903 ( .A(n1545), .B(n1543), .Y(n1823) );
  CLKINVX1 U904 ( .A(n1851), .Y(n1812) );
  CLKINVX1 U905 ( .A(n1811), .Y(n1857) );
  CLKINVX1 U906 ( .A(n1816), .Y(n1760) );
  AOI2BB1X1 U907 ( .A0N(n1752), .A1N(n1834), .B0(n861), .Y(n860) );
  AO21X1 U908 ( .A0(N71), .A1(n1868), .B0(n1751), .Y(n861) );
  AOI2BB1X1 U909 ( .A0N(n1789), .A1N(n1834), .B0(n863), .Y(n862) );
  AO21X1 U910 ( .A0(N69), .A1(n1868), .B0(n1788), .Y(n863) );
  AOI21XL U911 ( .A0(n128), .A1(n1836), .B0(n865), .Y(n864) );
  AO21X1 U912 ( .A0(N72), .A1(n1868), .B0(n1733), .Y(n865) );
  AOI21XL U913 ( .A0(n128), .A1(n1838), .B0(n867), .Y(n866) );
  AO21X1 U914 ( .A0(N70), .A1(n1868), .B0(n1771), .Y(n867) );
  NAND2XL U915 ( .A(n1348), .B(n1522), .Y(n1249) );
  NAND2XL U916 ( .A(N201), .B(n1515), .Y(n1247) );
  NAND3XL U917 ( .A(control[7]), .B(control[6]), .C(n1202), .Y(n1223) );
  NAND2X1 U918 ( .A(n1223), .B(n1222), .Y(n1464) );
  NAND2XL U919 ( .A(control[4]), .B(n1348), .Y(n1328) );
  MXI4X2 U920 ( .A(n1041), .B(n1042), .C(n1043), .D(n1044), .S0(N60), .S1(N59), 
        .Y(N105) );
  MXI4XL U921 ( .A(R4[10]), .B(R5[10]), .C(R6[10]), .D(R7[10]), .S0(N57), .S1(
        n1069), .Y(n1043) );
  MXI4XL U922 ( .A(R12[10]), .B(R13[10]), .C(R14[10]), .D(R15[10]), .S0(N57), 
        .S1(n1069), .Y(n1044) );
  MXI2X1 U923 ( .A(N104), .B(constant[11]), .S0(control[13]), .Y(n1350) );
  MXI4XL U924 ( .A(R4[11]), .B(R5[11]), .C(R6[11]), .D(R7[11]), .S0(N57), .S1(
        n1069), .Y(n1047) );
  MXI4XL U925 ( .A(R12[11]), .B(R13[11]), .C(R14[11]), .D(R15[11]), .S0(N57), 
        .S1(n1069), .Y(n1048) );
  MXI4XL U926 ( .A(R12[12]), .B(R13[12]), .C(R14[12]), .D(R15[12]), .S0(N57), 
        .S1(n1069), .Y(n1052) );
  MXI4XL U927 ( .A(R4[12]), .B(R5[12]), .C(R6[12]), .D(R7[12]), .S0(N57), .S1(
        n1069), .Y(n1051) );
  NAND2XL U928 ( .A(control[5]), .B(n1177), .Y(n1405) );
  NAND3X1 U929 ( .A(control[8]), .B(n1185), .C(n1221), .Y(n1484) );
  MXI4X1 U930 ( .A(R4[3]), .B(R5[3]), .C(R6[3]), .D(R7[3]), .S0(N57), .S1(
        n1066), .Y(n1015) );
  MXI4X1 U931 ( .A(R12[3]), .B(R13[3]), .C(R14[3]), .D(R15[3]), .S0(N57), .S1(
        n1066), .Y(n1016) );
  NAND3XL U932 ( .A(control[5]), .B(n1464), .C(n1462), .Y(n1313) );
  NAND2XL U933 ( .A(control[5]), .B(n1330), .Y(n1485) );
  MXI4X1 U934 ( .A(R12[4]), .B(R13[4]), .C(R14[4]), .D(R15[4]), .S0(N57), .S1(
        n1067), .Y(n1020) );
  MXI4X1 U935 ( .A(R4[4]), .B(R5[4]), .C(R6[4]), .D(R7[4]), .S0(N57), .S1(
        n1067), .Y(n1019) );
  MXI4XL U936 ( .A(R4[8]), .B(R5[8]), .C(R6[8]), .D(R7[8]), .S0(N57), .S1(
        n1068), .Y(n1035) );
  MXI4XL U937 ( .A(R12[8]), .B(R13[8]), .C(R14[8]), .D(R15[8]), .S0(N57), .S1(
        n1068), .Y(n1036) );
  AOI22XL U938 ( .A0(control[7]), .A1(n1186), .B0(control[8]), .B1(control[6]), 
        .Y(n869) );
  MXI4XL U939 ( .A(R8[15]), .B(R9[15]), .C(R10[15]), .D(R11[15]), .S0(N57), 
        .S1(n1070), .Y(n1062) );
  MXI4XL U940 ( .A(R12[15]), .B(R13[15]), .C(R14[15]), .D(R15[15]), .S0(N57), 
        .S1(n1070), .Y(n1064) );
  MXI4XL U941 ( .A(R0[15]), .B(R1[15]), .C(R2[15]), .D(R3[15]), .S0(N57), .S1(
        n1070), .Y(n1061) );
  CLKINVX1 U942 ( .A(control[5]), .Y(n1463) );
  MXI4X1 U943 ( .A(R8[1]), .B(R9[1]), .C(R10[1]), .D(R11[1]), .S0(n1138), .S1(
        n1146), .Y(n1078) );
  AND2XL U944 ( .A(n1482), .B(control[5]), .Y(n1489) );
  NAND2X1 U945 ( .A(control[3]), .B(n1175), .Y(n873) );
  NAND2XL U946 ( .A(N201), .B(control[3]), .Y(n874) );
  CLKBUFX3 U947 ( .A(N61), .Y(n1143) );
  NAND2X1 U948 ( .A(control[5]), .B(control[4]), .Y(n1530) );
  MXI2X1 U949 ( .A(n1549), .B(n919), .S0(control[11]), .Y(n1757) );
  NAND3X1 U950 ( .A(control[12]), .B(n1551), .C(n1550), .Y(n1816) );
  NAND2X1 U951 ( .A(n1545), .B(control[9]), .Y(n1795) );
  CLKINVX1 U952 ( .A(control[0]), .Y(n1868) );
  NOR2X1 U953 ( .A(N53), .B(N54), .Y(n90) );
  NOR2X1 U954 ( .A(n1176), .B(N54), .Y(n87) );
  NOR2BX1 U955 ( .AN(N54), .B(n1176), .Y(n94) );
  NOR2BX1 U956 ( .AN(N54), .B(N53), .Y(n97) );
  NOR2X1 U957 ( .A(n1866), .B(N55), .Y(n86) );
  NOR2X1 U958 ( .A(n1867), .B(N56), .Y(n93) );
  NOR2X1 U959 ( .A(N55), .B(N56), .Y(n105) );
  CLKINVX1 U960 ( .A(N53), .Y(n1176) );
  INVXL U961 ( .A(BUSB[1]), .Y(n1568) );
  NAND2XL U962 ( .A(n1759), .B(BUSB[1]), .Y(n1566) );
  CLKINVX1 U963 ( .A(BUSB[14]), .Y(n1802) );
  CLKINVX1 U964 ( .A(BUSB[5]), .Y(n1640) );
  CLKINVX1 U965 ( .A(BUSB[10]), .Y(n1722) );
  CLKINVX1 U966 ( .A(n1721), .Y(n1708) );
  CLKINVX1 U967 ( .A(BUSB[11]), .Y(n1741) );
  CLKINVX1 U968 ( .A(BUSB[2]), .Y(n1584) );
  CLKINVX1 U969 ( .A(BUSB[6]), .Y(n1657) );
  AND2X2 U970 ( .A(n1173), .B(n1815), .Y(n875) );
  CLKINVX1 U971 ( .A(n54), .Y(n1844) );
  NOR2X1 U972 ( .A(n1529), .B(n1528), .Y(n1532) );
  CLKINVX1 U973 ( .A(BUSB[13]), .Y(n1779) );
  CLKINVX1 U974 ( .A(BUSB[15]), .Y(n1817) );
  NAND2X1 U975 ( .A(n1759), .B(BUSB[5]), .Y(n1638) );
  NAND2X1 U976 ( .A(n1759), .B(BUSB[2]), .Y(n1582) );
  NAND2X1 U977 ( .A(n1759), .B(BUSB[6]), .Y(n1655) );
  CLKBUFX3 U978 ( .A(n992), .Y(n989) );
  CLKBUFX3 U979 ( .A(n992), .Y(n990) );
  CLKBUFX3 U980 ( .A(n991), .Y(n986) );
  CLKBUFX3 U981 ( .A(n991), .Y(n987) );
  CLKBUFX3 U982 ( .A(n992), .Y(n988) );
  CLKBUFX3 U983 ( .A(n991), .Y(n985) );
  NOR2X1 U984 ( .A(n1519), .B(n1518), .Y(n1535) );
  NAND4X1 U985 ( .A(n1414), .B(n1413), .C(n1412), .D(n1411), .Y(BUSB[7]) );
  AOI21X1 U986 ( .A0(n1499), .A1(n1498), .B0(n1497), .Y(n1510) );
  NOR3BXL U987 ( .AN(n1508), .B(n1507), .C(n1506), .Y(n1509) );
  NAND2X1 U988 ( .A(N209), .B(n1513), .Y(n1512) );
  NAND4X1 U989 ( .A(n1361), .B(n842), .C(n1360), .D(n1359), .Y(BUSB[10]) );
  NOR3X1 U990 ( .A(n1358), .B(n1357), .C(n1356), .Y(n1359) );
  AOI21X1 U991 ( .A0(N304), .A1(n1514), .B0(n1344), .Y(n1360) );
  AOI21X1 U992 ( .A0(N213), .A1(n1513), .B0(n1429), .Y(n1433) );
  NAND2X1 U993 ( .A(n1448), .B(n1447), .Y(n1453) );
  NAND4X1 U994 ( .A(n1394), .B(n841), .C(n1393), .D(n1392), .Y(BUSB[8]) );
  NAND2X1 U995 ( .A(n1238), .B(n1456), .Y(n1475) );
  NAND3X1 U996 ( .A(n1271), .B(n1270), .C(n1269), .Y(BUSB[14]) );
  NOR3X1 U997 ( .A(n1268), .B(n1267), .C(n1336), .Y(n1269) );
  AOI21X1 U998 ( .A0(N308), .A1(n1514), .B0(n1233), .Y(n1271) );
  NAND2X1 U999 ( .A(N221), .B(n1513), .Y(n1270) );
  NAND4X1 U1000 ( .A(n1380), .B(n843), .C(n1379), .D(n1378), .Y(BUSB[9]) );
  NOR4X1 U1001 ( .A(n1377), .B(n1376), .C(n1375), .D(n1374), .Y(n1378) );
  NAND4X1 U1002 ( .A(n1343), .B(n1342), .C(n1341), .D(n1340), .Y(BUSB[11]) );
  NOR2X1 U1003 ( .A(n1337), .B(n1336), .Y(n1342) );
  NOR2X1 U1004 ( .A(n1333), .B(n1332), .Y(n1343) );
  AOI22X1 U1005 ( .A0(n1338), .A1(n1498), .B0(N305), .B1(n1514), .Y(n1341) );
  NAND2X1 U1006 ( .A(n1383), .B(n1456), .Y(n1526) );
  NOR4X1 U1007 ( .A(n48), .B(n51), .C(n50), .D(n49), .Y(n1842) );
  AOI22X1 U1008 ( .A0(N298), .A1(n1514), .B0(n1448), .B1(n1466), .Y(n1467) );
  OAI2BB1X1 U1009 ( .A0N(N454), .A1N(n1857), .B0(n1579), .Y(n1591) );
  NAND2X1 U1010 ( .A(N435), .B(n900), .Y(n1579) );
  OAI2BB1X1 U1011 ( .A0N(N458), .A1N(n1857), .B0(n1652), .Y(n1664) );
  NAND2X1 U1012 ( .A(N439), .B(n900), .Y(n1652) );
  NOR2X1 U1013 ( .A(n1517), .B(n1430), .Y(n1431) );
  AOI22X1 U1014 ( .A0(N219), .A1(n1513), .B0(N306), .B1(n1514), .Y(n1318) );
  NOR3X1 U1015 ( .A(n1173), .B(n900), .C(n1859), .Y(n1864) );
  MXI2X1 U1016 ( .A(n899), .B(n1858), .S0(n892), .Y(n1859) );
  CLKINVX1 U1017 ( .A(BUSB[3]), .Y(n1602) );
  CLKINVX1 U1018 ( .A(BUSB[12]), .Y(n1758) );
  NAND3X1 U1019 ( .A(n1613), .B(n1612), .C(n1611), .Y(n49) );
  NOR2X1 U1020 ( .A(n1610), .B(n1609), .Y(n1611) );
  NAND2X1 U1021 ( .A(N555), .B(n1812), .Y(n1612) );
  AOI21X1 U1022 ( .A0(N516), .A1(n1852), .B0(n1595), .Y(n1613) );
  NAND3X1 U1023 ( .A(n1632), .B(n1631), .C(n1630), .Y(n50) );
  NOR2X1 U1024 ( .A(n1629), .B(n1628), .Y(n1630) );
  NAND2X1 U1025 ( .A(N556), .B(n1812), .Y(n1631) );
  AOI21X1 U1026 ( .A0(N517), .A1(n1852), .B0(n1614), .Y(n1632) );
  NAND3X1 U1027 ( .A(n1651), .B(n1650), .C(n1649), .Y(n51) );
  NOR2X1 U1028 ( .A(n1648), .B(n1647), .Y(n1649) );
  NAND2X1 U1029 ( .A(N557), .B(n1812), .Y(n1650) );
  AOI21X1 U1030 ( .A0(N518), .A1(n1852), .B0(n1633), .Y(n1651) );
  AOI21X1 U1031 ( .A0(N297), .A1(n1514), .B0(n1492), .Y(n1493) );
  AND2X2 U1032 ( .A(n1856), .B(n1568), .Y(n880) );
  AND2X2 U1033 ( .A(n1856), .B(n1621), .Y(n881) );
  AND2X2 U1034 ( .A(n1856), .B(n1758), .Y(n882) );
  AND2X2 U1035 ( .A(n1856), .B(n1689), .Y(n883) );
  AND2X2 U1036 ( .A(n1856), .B(n1722), .Y(n884) );
  AND2X2 U1037 ( .A(n1856), .B(n1741), .Y(n885) );
  AND2X2 U1038 ( .A(n1856), .B(n1802), .Y(n886) );
  AND2X2 U1039 ( .A(n1856), .B(n1673), .Y(n887) );
  AND2X2 U1040 ( .A(n1856), .B(n1707), .Y(n888) );
  AND2X2 U1041 ( .A(n1856), .B(n1552), .Y(n889) );
  NAND3X1 U1042 ( .A(n1731), .B(n1730), .C(n1729), .Y(n1836) );
  NAND2X1 U1043 ( .A(N562), .B(n1812), .Y(n1730) );
  AOI21X1 U1044 ( .A0(N523), .A1(n1852), .B0(n1718), .Y(n1731) );
  NOR2X1 U1045 ( .A(n1728), .B(n1727), .Y(n1729) );
  NAND3X1 U1046 ( .A(n1769), .B(n1768), .C(n1767), .Y(n1838) );
  AOI21X1 U1047 ( .A0(N525), .A1(n1852), .B0(n1753), .Y(n1769) );
  NAND2X1 U1048 ( .A(N564), .B(n1812), .Y(n1768) );
  NOR2X1 U1049 ( .A(n1766), .B(n1765), .Y(n1767) );
  NAND3X1 U1050 ( .A(n1699), .B(n1698), .C(n1697), .Y(n54) );
  NAND2X1 U1051 ( .A(N560), .B(n1812), .Y(n1698) );
  AOI21X1 U1052 ( .A0(N521), .A1(n1852), .B0(n1684), .Y(n1699) );
  NOR2X1 U1053 ( .A(n1696), .B(n1695), .Y(n1697) );
  NAND2X1 U1054 ( .A(N217), .B(n1513), .Y(n1361) );
  NAND3X1 U1055 ( .A(n1807), .B(n1806), .C(n1805), .Y(n1840) );
  AOI21X1 U1056 ( .A0(N527), .A1(n1852), .B0(n1790), .Y(n1807) );
  AOI21X1 U1057 ( .A0(N566), .A1(n1812), .B0(n1796), .Y(n1806) );
  NOR4X1 U1058 ( .A(n1804), .B(n894), .C(n875), .D(n1803), .Y(n1805) );
  OAI2BB1X1 U1059 ( .A0N(N464), .A1N(n1857), .B0(n1754), .Y(n1766) );
  NAND2X1 U1060 ( .A(N445), .B(n900), .Y(n1754) );
  OAI2BB1X1 U1061 ( .A0N(N459), .A1N(n1857), .B0(n1668), .Y(n1680) );
  NAND2X1 U1062 ( .A(N440), .B(n900), .Y(n1668) );
  OAI2BB1X1 U1063 ( .A0N(N462), .A1N(n1857), .B0(n1719), .Y(n1728) );
  NAND2X1 U1064 ( .A(N443), .B(n900), .Y(n1719) );
  NOR2X1 U1065 ( .A(n53), .B(n52), .Y(n1843) );
  NAND2X1 U1066 ( .A(n1686), .B(n1685), .Y(n1696) );
  NAND2X1 U1067 ( .A(N441), .B(n900), .Y(n1685) );
  NAND2X1 U1068 ( .A(N460), .B(n1857), .Y(n1686) );
  NAND2X1 U1069 ( .A(n1597), .B(n1596), .Y(n1610) );
  NAND2X1 U1070 ( .A(N436), .B(n900), .Y(n1596) );
  NAND2X1 U1071 ( .A(N455), .B(n1857), .Y(n1597) );
  NAND2X1 U1072 ( .A(n1616), .B(n1615), .Y(n1629) );
  NAND2X1 U1073 ( .A(N437), .B(n900), .Y(n1615) );
  NAND2X1 U1074 ( .A(N456), .B(n1857), .Y(n1616) );
  NAND2X1 U1075 ( .A(n1635), .B(n1634), .Y(n1648) );
  NAND2X1 U1076 ( .A(N438), .B(n900), .Y(n1634) );
  NAND2X1 U1077 ( .A(N457), .B(n1857), .Y(n1635) );
  CLKINVX1 U1078 ( .A(n1178), .Y(n1177) );
  CLKBUFX3 U1079 ( .A(n1444), .Y(n1162) );
  NAND2X1 U1080 ( .A(n1173), .B(n1669), .Y(n1670) );
  CLKINVX1 U1081 ( .A(\add_233/carry[7] ), .Y(n1669) );
  CLKINVX1 U1082 ( .A(n1791), .Y(n1798) );
  AND2X2 U1083 ( .A(N502), .B(n901), .Y(n1746) );
  AND2X2 U1084 ( .A(N500), .B(n901), .Y(n1710) );
  CLKINVX1 U1085 ( .A(\FUResult[15] ), .Y(n1862) );
  NAND2X1 U1086 ( .A(N294), .B(n1514), .Y(n1205) );
  NAND2X1 U1087 ( .A(N507), .B(n901), .Y(n1850) );
  CLKINVX1 U1088 ( .A(n1186), .Y(n1202) );
  MXI2X1 U1089 ( .A(n1760), .B(n1759), .S0(n1689), .Y(n1690) );
  MXI2X1 U1090 ( .A(n1760), .B(n1759), .S0(n1722), .Y(n1723) );
  MXI2X1 U1091 ( .A(n1760), .B(n1759), .S0(n1758), .Y(n1761) );
  CLKINVX1 U1092 ( .A(n1847), .Y(n1815) );
  AND2X2 U1093 ( .A(N506), .B(n901), .Y(n1826) );
  CLKINVX1 U1094 ( .A(n1483), .Y(n1488) );
  OAI2BB1X1 U1095 ( .A0N(N453), .A1N(n1857), .B0(n1564), .Y(n1575) );
  NAND2XL U1096 ( .A(N434), .B(n900), .Y(n1564) );
  NOR2BX1 U1097 ( .AN(n1846), .B(n1845), .Y(Z) );
  NOR4BX1 U1098 ( .AN(n1841), .B(n1840), .C(n839), .D(n1839), .Y(n1846) );
  NAND4X1 U1099 ( .A(n1844), .B(n1862), .C(n1843), .D(n1842), .Y(n1845) );
  NOR4X1 U1100 ( .A(n1836), .B(n1835), .C(n47), .D(n41), .Y(n1841) );
  CLKINVX1 U1101 ( .A(N463), .Y(n1734) );
  CLKINVX1 U1102 ( .A(N461), .Y(n1700) );
  CLKINVX1 U1103 ( .A(N465), .Y(n1772) );
  CLKINVX1 U1104 ( .A(n1472), .Y(n1473) );
  NAND3X1 U1105 ( .A(n1232), .B(n1231), .C(n1230), .Y(BUSB[15]) );
  NOR3X1 U1106 ( .A(n1229), .B(n1228), .C(n1227), .Y(n1230) );
  NAND2X1 U1107 ( .A(N309), .B(n1514), .Y(n1231) );
  NAND2X1 U1108 ( .A(N222), .B(n1513), .Y(n1232) );
  NAND3X1 U1109 ( .A(n1299), .B(n1298), .C(n1297), .Y(BUSB[13]) );
  NOR3X1 U1110 ( .A(n1296), .B(n1295), .C(n1336), .Y(n1297) );
  AOI21X1 U1111 ( .A0(N307), .A1(n1514), .B0(n1272), .Y(n1299) );
  NAND2X1 U1112 ( .A(N220), .B(n1513), .Y(n1298) );
  OAI22XL U1113 ( .A0(n856), .A1(n1335), .B0(n1282), .B1(n1517), .Y(n1296) );
  OAI22XL U1114 ( .A0(n1395), .A1(n1435), .B0(n1491), .B1(n1373), .Y(n1333) );
  OAI22XL U1115 ( .A0(n1355), .A1(n1517), .B0(n1475), .B1(n1505), .Y(n1358) );
  CLKINVX1 U1116 ( .A(n1345), .Y(n1355) );
  OAI22XL U1117 ( .A0(n1404), .A1(n1475), .B0(n1491), .B1(n1435), .Y(n1410) );
  CLKINVX1 U1118 ( .A(n1478), .Y(n1404) );
  NAND4X1 U1119 ( .A(n1563), .B(n1562), .C(n1561), .D(n1560), .Y(n41) );
  NAND2X1 U1120 ( .A(N552), .B(n1812), .Y(n1561) );
  NAND2X1 U1121 ( .A(N513), .B(n1852), .Y(n1562) );
  CLKINVX1 U1122 ( .A(n857), .Y(n1423) );
  AND2X2 U1123 ( .A(n1856), .B(n1779), .Y(n890) );
  AND2X2 U1124 ( .A(n1856), .B(n1817), .Y(n891) );
  CLKINVX1 U1125 ( .A(n1517), .Y(n1498) );
  NAND2X1 U1126 ( .A(n1759), .B(BUSB[3]), .Y(n1600) );
  NOR2BX1 U1127 ( .AN(n1370), .B(n1517), .Y(n1376) );
  NAND2X1 U1128 ( .A(n1457), .B(n1456), .Y(n1528) );
  NOR2X1 U1129 ( .A(n892), .B(n1823), .Y(n1824) );
  NAND2X1 U1130 ( .A(n1369), .B(n1368), .Y(n1434) );
  NAND2X1 U1131 ( .A(n1198), .B(n1197), .Y(n1388) );
  NAND2X1 U1132 ( .A(n1291), .B(n1290), .Y(n1370) );
  NOR2X1 U1133 ( .A(n1401), .B(n1472), .Y(n1290) );
  NOR2X1 U1134 ( .A(n1365), .B(n1442), .Y(n1291) );
  CLKINVX1 U1135 ( .A(n1335), .Y(n1238) );
  NAND2X1 U1136 ( .A(n1220), .B(n1219), .Y(n1338) );
  NOR2X1 U1137 ( .A(n1322), .B(n1399), .Y(n1220) );
  NOR2X1 U1138 ( .A(n1367), .B(n1439), .Y(n1219) );
  NOR2X1 U1139 ( .A(n1559), .B(n1558), .Y(n1560) );
  NAND2X1 U1140 ( .A(n1541), .B(n1540), .Y(n1559) );
  NAND2X1 U1141 ( .A(n1557), .B(n1556), .Y(n1558) );
  NAND2XL U1142 ( .A(N433), .B(n900), .Y(n1540) );
  NOR2X1 U1143 ( .A(n1505), .B(n1528), .Y(n1506) );
  NAND2XL U1144 ( .A(N449), .B(n900), .Y(n1848) );
  NAND2X1 U1145 ( .A(n1173), .B(n1617), .Y(n1618) );
  CLKINVX1 U1146 ( .A(\add_233/carry[4] ), .Y(n1617) );
  NAND2X1 U1147 ( .A(n1173), .B(n1653), .Y(n1654) );
  CLKINVX1 U1148 ( .A(\add_233/carry[6] ), .Y(n1653) );
  NAND2X1 U1149 ( .A(n1246), .B(n1245), .Y(n1268) );
  NAND2X1 U1150 ( .A(n1243), .B(n1242), .Y(n1244) );
  NAND2X1 U1151 ( .A(N452), .B(n1857), .Y(n1541) );
  XOR2X1 U1152 ( .A(BUSB[15]), .B(n1861), .Y(n892) );
  CLKBUFX3 U1153 ( .A(n1444), .Y(n1163) );
  CLKINVX1 U1154 ( .A(n1371), .Y(n1450) );
  CLKINVX1 U1155 ( .A(n1395), .Y(n1396) );
  AND2X2 U1156 ( .A(N444), .B(n900), .Y(n893) );
  AND2X2 U1157 ( .A(N447), .B(n900), .Y(n894) );
  AND2X2 U1158 ( .A(N446), .B(n900), .Y(n895) );
  AND2X2 U1159 ( .A(N442), .B(n900), .Y(n896) );
  AND2X2 U1160 ( .A(N448), .B(n900), .Y(n897) );
  NAND2X1 U1161 ( .A(n1173), .B(n1636), .Y(n1637) );
  CLKINVX1 U1162 ( .A(\add_233/carry[5] ), .Y(n1636) );
  NOR2BX1 U1163 ( .AN(n1381), .B(n1517), .Y(n1382) );
  CLKINVX1 U1164 ( .A(n1527), .Y(n1447) );
  NOR2X1 U1165 ( .A(n1226), .B(n1517), .Y(n1227) );
  NAND2X1 U1166 ( .A(n1174), .B(n1598), .Y(n1599) );
  CLKINVX1 U1167 ( .A(\add_233/carry[3] ), .Y(n1598) );
  CLKINVX1 U1168 ( .A(n1547), .Y(n1544) );
  NAND2X1 U1169 ( .A(n1174), .B(n1580), .Y(n1581) );
  CLKINVX1 U1170 ( .A(\add_233/carry[2] ), .Y(n1580) );
  CLKBUFX3 U1171 ( .A(n1860), .Y(n1173) );
  CLKBUFX3 U1172 ( .A(n1860), .Y(n1174) );
  NOR2X1 U1173 ( .A(n901), .B(n1857), .Y(n1858) );
  CLKBUFX3 U1174 ( .A(N53), .Y(n992) );
  CLKBUFX3 U1175 ( .A(N53), .Y(n991) );
  OAI21XL U1176 ( .A0(n1744), .A1(n1814), .B0(n1757), .Y(n1735) );
  NOR2X1 U1177 ( .A(n1780), .B(n1814), .Y(n1755) );
  NAND3BX1 U1178 ( .AN(n1481), .B(n1480), .C(n1479), .Y(n1495) );
  AOI21X1 U1179 ( .A0(N210), .A1(n1513), .B0(n1490), .Y(n1494) );
  AOI22X1 U1180 ( .A0(n1317), .A1(MUXB[12]), .B0(n1448), .B1(n1316), .Y(n1319)
         );
  NAND3X1 U1181 ( .A(n1315), .B(n1314), .C(n1313), .Y(n1320) );
  NOR2X1 U1182 ( .A(n1791), .B(n1814), .Y(n1781) );
  NOR2X1 U1183 ( .A(n1406), .B(n1328), .Y(n1329) );
  NOR3X1 U1184 ( .A(n1490), .B(n1461), .C(n1460), .Y(n1470) );
  NAND3X1 U1185 ( .A(n1464), .B(n1463), .C(n1462), .Y(n1469) );
  AOI21X1 U1186 ( .A0(N211), .A1(n1513), .B0(n1465), .Y(n1468) );
  CLKINVX1 U1187 ( .A(BUSA[10]), .Y(n1743) );
  CLKINVX1 U1188 ( .A(BUSA[11]), .Y(n1742) );
  NAND3X1 U1189 ( .A(n1185), .B(n1221), .C(n1183), .Y(n1184) );
  NAND4BX2 U1190 ( .AN(n1207), .B(n1206), .C(n1205), .D(n1204), .Y(BUSB[0]) );
  OAI22XL U1191 ( .A0(n1187), .A1(n1475), .B0(n1384), .B1(n898), .Y(n1207) );
  OAI21XL U1192 ( .A0(n1201), .A1(n1200), .B0(n1456), .Y(n1206) );
  NAND2X1 U1193 ( .A(N207), .B(n1513), .Y(n1204) );
  OAI2BB1X1 U1194 ( .A0N(N493), .A1N(n901), .B0(n1589), .Y(n1590) );
  MXI2X1 U1195 ( .A(n1588), .B(n1587), .S0(BUSA[2]), .Y(n1589) );
  NAND3X1 U1196 ( .A(n1582), .B(n1795), .C(n1581), .Y(n1588) );
  OAI2BB1X1 U1197 ( .A0N(N497), .A1N(n901), .B0(n1662), .Y(n1663) );
  MXI2X1 U1198 ( .A(n1661), .B(n1660), .S0(BUSA[6]), .Y(n1662) );
  NAND3X1 U1199 ( .A(n1655), .B(n1795), .C(n1654), .Y(n1661) );
  NAND4X1 U1200 ( .A(n1212), .B(n1211), .C(n1210), .D(n1209), .Y(n1491) );
  OR2X1 U1201 ( .A(BUSA[5]), .B(\add_233/carry[5] ), .Y(\add_233/carry[6] ) );
  MXI2X1 U1202 ( .A(n1822), .B(n1821), .S0(BUSA[15]), .Y(n1825) );
  NOR3X1 U1203 ( .A(n1820), .B(n1819), .C(n1818), .Y(n1821) );
  NOR2X1 U1204 ( .A(n1813), .B(n875), .Y(n1822) );
  NOR2X1 U1205 ( .A(n1817), .B(n1816), .Y(n1818) );
  AOI21X1 U1206 ( .A0(N218), .A1(n1513), .B0(n1339), .Y(n1340) );
  NOR2X1 U1207 ( .A(n1350), .B(n869), .Y(n1339) );
  NOR3X1 U1208 ( .A(\add_233/carry[8] ), .B(BUSA[9]), .C(BUSA[8]), .Y(n1744)
         );
  OAI21XL U1209 ( .A0(n1527), .A1(n1526), .B0(n1525), .Y(n1533) );
  OAI21XL U1210 ( .A0(n1524), .A1(n1523), .B0(n1448), .Y(n1525) );
  OAI22XL U1211 ( .A0(n1522), .A1(n857), .B0(n1521), .B1(n873), .Y(n1523) );
  NAND2X1 U1212 ( .A(n1694), .B(n1693), .Y(n1695) );
  NAND2X1 U1213 ( .A(N499), .B(n901), .Y(n1694) );
  MXI2X1 U1214 ( .A(n1692), .B(n1691), .S0(BUSA[8]), .Y(n1693) );
  NAND2X1 U1215 ( .A(n1163), .B(n1330), .Y(n1179) );
  MXI2X1 U1216 ( .A(n1795), .B(n1737), .S0(BUSA[11]), .Y(n1738) );
  NOR3X1 U1217 ( .A(n1736), .B(n844), .C(n1735), .Y(n1737) );
  MXI2X1 U1218 ( .A(n1816), .B(n1823), .S0(n1741), .Y(n1736) );
  MXI2X1 U1219 ( .A(n1795), .B(n1794), .S0(BUSA[14]), .Y(n1796) );
  NOR3X1 U1220 ( .A(n1793), .B(n1792), .C(n1820), .Y(n1794) );
  MXI2X1 U1221 ( .A(n1816), .B(n1823), .S0(n1802), .Y(n1793) );
  NOR2X1 U1222 ( .A(n1798), .B(n1814), .Y(n1792) );
  NAND4X1 U1223 ( .A(n1279), .B(n1278), .C(n1277), .D(n1276), .Y(n1280) );
  NOR3X1 U1224 ( .A(n1275), .B(n1274), .C(n1273), .Y(n1281) );
  OAI2BB1X1 U1225 ( .A0N(n1174), .A1N(n1780), .B0(n1757), .Y(n1773) );
  OAI21XL U1226 ( .A0(BUSA[15]), .A1(n1847), .B0(n1174), .Y(n1849) );
  NAND2BX1 U1227 ( .AN(n1570), .B(n1569), .Y(n1571) );
  NAND2X1 U1228 ( .A(n1757), .B(n1567), .Y(n1570) );
  MXI2X1 U1229 ( .A(n1760), .B(n1759), .S0(n1568), .Y(n1569) );
  NAND2X1 U1230 ( .A(BUSA[0]), .B(n1173), .Y(n1567) );
  NAND3X1 U1231 ( .A(n1713), .B(n1712), .C(n1711), .Y(n1835) );
  AOI2BB2X1 U1232 ( .B0(N522), .B1(n1852), .A0N(n1811), .A1N(n1700), .Y(n1713)
         );
  AOI21X1 U1233 ( .A0(N561), .A1(n1812), .B0(n1704), .Y(n1712) );
  NOR4X1 U1234 ( .A(n1710), .B(n896), .C(n1709), .D(n1708), .Y(n1711) );
  NAND3X1 U1235 ( .A(n1594), .B(n1593), .C(n1592), .Y(n48) );
  NOR2X1 U1236 ( .A(n1591), .B(n1590), .Y(n1592) );
  NAND2BX1 U1237 ( .AN(n1851), .B(N554), .Y(n1593) );
  NAND3X1 U1238 ( .A(n1578), .B(n1577), .C(n1576), .Y(n47) );
  NOR2X1 U1239 ( .A(n1575), .B(n1574), .Y(n1576) );
  NAND2BX1 U1240 ( .AN(n1851), .B(N553), .Y(n1577) );
  AOI2BB2X1 U1241 ( .B0(N514), .B1(n1852), .A0N(n1568), .A1N(n847), .Y(n1578)
         );
  NAND3X1 U1242 ( .A(n1667), .B(n1666), .C(n1665), .Y(n52) );
  NOR2X1 U1243 ( .A(n1664), .B(n1663), .Y(n1665) );
  NAND2BX1 U1244 ( .AN(n1851), .B(N558), .Y(n1666) );
  NAND3X1 U1245 ( .A(n1683), .B(n1682), .C(n1681), .Y(n53) );
  NOR2X1 U1246 ( .A(n1680), .B(n1679), .Y(n1681) );
  NAND2BX1 U1247 ( .AN(n1851), .B(N559), .Y(n1682) );
  NAND2X1 U1248 ( .A(n1177), .B(n1463), .Y(n1471) );
  OAI21XL U1249 ( .A0(n1526), .A1(n1504), .B0(n1503), .Y(n1507) );
  OAI21XL U1250 ( .A0(n1502), .A1(n1501), .B0(n1448), .Y(n1503) );
  OAI22XL U1251 ( .A0(n1521), .A1(n857), .B0(n1520), .B1(n873), .Y(n1501) );
  NAND2BX1 U1252 ( .AN(n1675), .B(n1674), .Y(n1676) );
  NAND2X1 U1253 ( .A(n1757), .B(n1672), .Y(n1675) );
  NAND2X1 U1254 ( .A(\add_233/carry[7] ), .B(n1173), .Y(n1672) );
  NAND2X1 U1255 ( .A(n873), .B(n857), .Y(N202) );
  NAND3X1 U1256 ( .A(n1749), .B(n1748), .C(n1747), .Y(n1837) );
  AOI2BB2X1 U1257 ( .B0(N524), .B1(n1852), .A0N(n1811), .A1N(n1734), .Y(n1749)
         );
  NOR4X1 U1258 ( .A(n1746), .B(n893), .C(n1745), .D(n1755), .Y(n1747) );
  AOI21X1 U1259 ( .A0(N563), .A1(n1812), .B0(n1738), .Y(n1748) );
  NAND3X1 U1260 ( .A(n1721), .B(n1795), .C(n1720), .Y(n1725) );
  NAND2X1 U1261 ( .A(n1759), .B(BUSB[10]), .Y(n1720) );
  NAND2X1 U1262 ( .A(n1237), .B(n1236), .Y(n1500) );
  NAND2X1 U1263 ( .A(n1264), .B(n1235), .Y(n1236) );
  NAND2X1 U1264 ( .A(n1757), .B(n1688), .Y(n1701) );
  NAND2X1 U1265 ( .A(\add_233/carry[8] ), .B(n1173), .Y(n1688) );
  OAI21XL U1266 ( .A0(n1477), .A1(n1476), .B0(n1448), .Y(n1480) );
  NOR2XL U1267 ( .A(n1520), .B(n857), .Y(n1477) );
  OAI21XL U1268 ( .A0(n1474), .A1(n873), .B0(n1473), .Y(n1476) );
  NOR2X1 U1269 ( .A(n1346), .B(n857), .Y(n1325) );
  NAND3X1 U1270 ( .A(n1786), .B(n1785), .C(n1784), .Y(n1839) );
  AOI2BB2X1 U1271 ( .B0(N526), .B1(n1852), .A0N(n1811), .A1N(n1772), .Y(n1786)
         );
  NOR4X1 U1272 ( .A(n1783), .B(n895), .C(n1782), .D(n1781), .Y(n1784) );
  AOI21X1 U1273 ( .A0(N565), .A1(n1812), .B0(n1776), .Y(n1785) );
  NOR2X1 U1274 ( .A(n856), .B(n1530), .Y(n1531) );
  NOR3X1 U1275 ( .A(n1486), .B(n1485), .C(n1484), .Y(n1487) );
  NOR2XL U1276 ( .A(n1420), .B(n873), .Y(n1399) );
  NOR2X1 U1277 ( .A(n1418), .B(n857), .Y(n1401) );
  NOR2X1 U1278 ( .A(n1815), .B(n1814), .Y(n1819) );
  NAND2X1 U1279 ( .A(n1403), .B(n1402), .Y(n1478) );
  NOR2X1 U1280 ( .A(n1422), .B(n1163), .Y(n1398) );
  MXI2X1 U1281 ( .A(n1795), .B(n1775), .S0(BUSA[13]), .Y(n1776) );
  NOR3X1 U1282 ( .A(n1774), .B(n845), .C(n1773), .Y(n1775) );
  MXI2X1 U1283 ( .A(n1816), .B(n1823), .S0(n1779), .Y(n1774) );
  AOI2BB2X1 U1284 ( .B0(N567), .B1(n1812), .A0N(n1817), .A1N(n847), .Y(n1828)
         );
  MXI2X1 U1285 ( .A(n1795), .B(n1703), .S0(BUSA[9]), .Y(n1704) );
  NOR3X1 U1286 ( .A(n1702), .B(n846), .C(n1701), .Y(n1703) );
  MXI2X1 U1287 ( .A(n1816), .B(n1823), .S0(n1707), .Y(n1702) );
  NAND2X1 U1288 ( .A(n1759), .B(BUSB[12]), .Y(n1756) );
  NAND2X1 U1289 ( .A(n1471), .B(n1183), .Y(n1186) );
  NAND2X1 U1290 ( .A(n1327), .B(n1326), .Y(n1334) );
  OAI2BB1X1 U1291 ( .A0N(N498), .A1N(n901), .B0(n1678), .Y(n1679) );
  MXI2X1 U1292 ( .A(n1677), .B(n1676), .S0(BUSA[7]), .Y(n1678) );
  NAND3X1 U1293 ( .A(n1671), .B(n1795), .C(n1670), .Y(n1677) );
  OAI2BB1X1 U1294 ( .A0N(N492), .A1N(n901), .B0(n1573), .Y(n1574) );
  MXI2X1 U1295 ( .A(n1572), .B(n1571), .S0(BUSA[1]), .Y(n1573) );
  NAND3X1 U1296 ( .A(n1566), .B(n1795), .C(n1565), .Y(n1572) );
  CLKINVX1 U1297 ( .A(n1372), .Y(n1415) );
  CLKINVX1 U1298 ( .A(BUSA[14]), .Y(n1797) );
  OAI2BB1X1 U1299 ( .A0N(N503), .A1N(n901), .B0(n1764), .Y(n1765) );
  MXI2X1 U1300 ( .A(n1763), .B(n1762), .S0(BUSA[12]), .Y(n1764) );
  OAI2BB1X1 U1301 ( .A0N(N501), .A1N(n901), .B0(n1726), .Y(n1727) );
  MXI2X1 U1302 ( .A(n1725), .B(n1724), .S0(BUSA[10]), .Y(n1726) );
  NAND2X1 U1303 ( .A(n1627), .B(n1626), .Y(n1628) );
  MXI2X1 U1304 ( .A(n1625), .B(n1624), .S0(BUSA[4]), .Y(n1626) );
  NAND2X1 U1305 ( .A(N495), .B(n901), .Y(n1627) );
  NAND3X1 U1306 ( .A(n1619), .B(n1795), .C(n1618), .Y(n1625) );
  NAND2X1 U1307 ( .A(n1646), .B(n1645), .Y(n1647) );
  MXI2X1 U1308 ( .A(n1644), .B(n1643), .S0(BUSA[5]), .Y(n1645) );
  NAND2X1 U1309 ( .A(N496), .B(n901), .Y(n1646) );
  NAND3X1 U1310 ( .A(n1638), .B(n1795), .C(n1637), .Y(n1644) );
  NAND2X1 U1311 ( .A(n1608), .B(n1607), .Y(n1609) );
  MXI2X1 U1312 ( .A(n1606), .B(n1605), .S0(BUSA[3]), .Y(n1607) );
  NAND2X1 U1313 ( .A(N494), .B(n901), .Y(n1608) );
  NAND3X1 U1314 ( .A(n1600), .B(n1795), .C(n1599), .Y(n1606) );
  CLKINVX1 U1315 ( .A(n1520), .Y(MUXB[4]) );
  CLKINVX1 U1316 ( .A(n1346), .Y(MUXB[12]) );
  NAND3BX1 U1317 ( .AN(n1855), .B(n1854), .C(n1853), .Y(C) );
  NAND3X1 U1318 ( .A(n1850), .B(n1849), .C(n1848), .Y(n1855) );
  AOI22X1 U1319 ( .A0(N468), .A1(n1857), .B0(N529), .B1(n1852), .Y(n1853) );
  NAND2BX1 U1320 ( .AN(n1851), .B(N568), .Y(n1854) );
  CLKBUFX3 U1321 ( .A(n1143), .Y(n1138) );
  NAND2X1 U1322 ( .A(n1348), .B(n1330), .Y(n1178) );
  CLKINVX1 U1323 ( .A(n1323), .Y(MUXB[14]) );
  CLKINVX1 U1324 ( .A(n1474), .Y(MUXB[5]) );
  CLKINVX1 U1325 ( .A(n1521), .Y(MUXB[3]) );
  CLKINVX1 U1326 ( .A(n1422), .Y(MUXB[7]) );
  CLKINVX1 U1327 ( .A(n1420), .Y(MUXB[9]) );
  CLKINVX1 U1328 ( .A(n1418), .Y(MUXB[8]) );
  NAND2BX1 U1329 ( .AN(n1530), .B(n1500), .Y(n1508) );
  CLKBUFX3 U1330 ( .A(n1071), .Y(n1067) );
  CLKBUFX3 U1331 ( .A(n1072), .Y(n1068) );
  CLKBUFX3 U1332 ( .A(n1072), .Y(n1070) );
  CLKBUFX3 U1333 ( .A(n1071), .Y(n1066) );
  CLKBUFX3 U1334 ( .A(n1072), .Y(n1069) );
  CLKBUFX3 U1335 ( .A(n1151), .Y(n1146) );
  CLKBUFX3 U1336 ( .A(n1143), .Y(n1137) );
  CLKBUFX3 U1337 ( .A(n1071), .Y(n1065) );
  CLKBUFX3 U1338 ( .A(n1151), .Y(n1145) );
  NAND4X1 U1339 ( .A(n1427), .B(n1426), .C(n1425), .D(n1424), .Y(n1504) );
  NAND2X1 U1340 ( .A(n1419), .B(n1418), .Y(n1427) );
  NAND2X1 U1341 ( .A(n1421), .B(n1420), .Y(n1425) );
  NAND2X1 U1342 ( .A(n1423), .B(n1422), .Y(n1424) );
  NAND4X1 U1343 ( .A(n1312), .B(n1311), .C(n1310), .D(n1309), .Y(n1387) );
  NAND2X1 U1344 ( .A(n1423), .B(n1521), .Y(n1309) );
  NAND4X1 U1345 ( .A(n1354), .B(n1353), .C(n1352), .D(n1351), .Y(n1505) );
  NAND2X1 U1346 ( .A(n1419), .B(n1346), .Y(n1354) );
  OAI21XL U1347 ( .A0(n1435), .A1(n1516), .B0(n1455), .Y(n1436) );
  NAND4X1 U1348 ( .A(n1216), .B(n1215), .C(n1214), .D(n1213), .Y(n1395) );
  NAND2X1 U1349 ( .A(n1419), .B(n1474), .Y(n1216) );
  AOI21X1 U1350 ( .A0(n1294), .A1(n1293), .B0(n1292), .Y(n1295) );
  NAND2X1 U1351 ( .A(n1383), .B(n1370), .Y(n1293) );
  AOI21X1 U1352 ( .A0(n1262), .A1(n1261), .B0(n1292), .Y(n1267) );
  NAND2X1 U1353 ( .A(n1383), .B(n1345), .Y(n1261) );
  NOR2X1 U1354 ( .A(n1254), .B(n1253), .Y(n1262) );
  AOI21X1 U1355 ( .A0(n1225), .A1(n1224), .B0(n1292), .Y(n1228) );
  NAND2X1 U1356 ( .A(n1383), .B(n1338), .Y(n1224) );
  NOR2X1 U1357 ( .A(n1218), .B(n1217), .Y(n1225) );
  MXI2X1 U1358 ( .A(n1555), .B(n1554), .S0(BUSA[0]), .Y(n1556) );
  OAI21XL U1359 ( .A0(n1552), .A1(n1823), .B0(n1546), .Y(n1555) );
  NAND2BX1 U1360 ( .AN(n1820), .B(n1553), .Y(n1554) );
  NOR2X1 U1361 ( .A(n1174), .B(n1813), .Y(n1546) );
  INVX1 U1362 ( .A(n874), .Y(n1421) );
  INVX1 U1363 ( .A(n873), .Y(n1419) );
  OAI21XL U1364 ( .A0(n1516), .A1(n1373), .B0(n1372), .Y(n1374) );
  OAI21XL U1365 ( .A0(n1458), .A1(n1526), .B0(n1386), .Y(n1391) );
  NAND2X1 U1366 ( .A(N491), .B(n901), .Y(n1557) );
  OAI21XL U1367 ( .A0(n1496), .A1(n1373), .B0(n1372), .Y(n1356) );
  NOR2X1 U1368 ( .A(n1406), .B(n1265), .Y(n1266) );
  NAND2X1 U1369 ( .A(n1264), .B(n1383), .Y(n1265) );
  NAND2X1 U1370 ( .A(n1288), .B(n1287), .Y(n1516) );
  NAND4X1 U1371 ( .A(n1286), .B(n1285), .C(n1284), .D(n1283), .Y(n1371) );
  NAND2X1 U1372 ( .A(n1419), .B(n1521), .Y(n1286) );
  NAND2BX1 U1373 ( .AN(n1586), .B(n1585), .Y(n1587) );
  NAND2X1 U1374 ( .A(n1757), .B(n1583), .Y(n1586) );
  NAND2X1 U1375 ( .A(\add_233/carry[2] ), .B(n1173), .Y(n1583) );
  NAND2BX1 U1376 ( .AN(n1604), .B(n1603), .Y(n1605) );
  NAND2X1 U1377 ( .A(n1757), .B(n1601), .Y(n1604) );
  NAND2X1 U1378 ( .A(\add_233/carry[3] ), .B(n1173), .Y(n1601) );
  NAND2BX1 U1379 ( .AN(n1623), .B(n1622), .Y(n1624) );
  NAND2X1 U1380 ( .A(n1757), .B(n1620), .Y(n1623) );
  NAND2X1 U1381 ( .A(\add_233/carry[4] ), .B(n1173), .Y(n1620) );
  NAND2BX1 U1382 ( .AN(n1642), .B(n1641), .Y(n1643) );
  NAND2X1 U1383 ( .A(n1757), .B(n1639), .Y(n1642) );
  NAND2X1 U1384 ( .A(\add_233/carry[5] ), .B(n1173), .Y(n1639) );
  NAND2BX1 U1385 ( .AN(n1659), .B(n1658), .Y(n1660) );
  NAND2X1 U1386 ( .A(n1757), .B(n1656), .Y(n1659) );
  OAI21XL U1387 ( .A0(n1303), .A1(n1302), .B0(n1498), .Y(n1315) );
  NOR2XL U1388 ( .A(n1420), .B(n874), .Y(n1303) );
  OAI21XL U1389 ( .A0(n1350), .A1(n857), .B0(n1301), .Y(n1302) );
  OAI21XL U1390 ( .A0(n1486), .A1(n1526), .B0(n1408), .Y(n1409) );
  NOR2X1 U1391 ( .A(n1406), .B(n1405), .Y(n1407) );
  NOR2X1 U1392 ( .A(n1422), .B(n873), .Y(n1442) );
  NOR2XL U1393 ( .A(n1418), .B(n874), .Y(n1439) );
  CLKINVX1 U1394 ( .A(n1484), .Y(n1264) );
  NOR2X1 U1395 ( .A(n1802), .B(n1801), .Y(n1803) );
  NOR2X1 U1396 ( .A(n1800), .B(n1799), .Y(n1801) );
  NOR2X1 U1397 ( .A(BUSA[14]), .B(n1823), .Y(n1799) );
  OAI21XL U1398 ( .A0(n1458), .A1(n1530), .B0(n1199), .Y(n1200) );
  NOR2X1 U1399 ( .A(n1741), .B(n1740), .Y(n1745) );
  NOR2X1 U1400 ( .A(n1800), .B(n1739), .Y(n1740) );
  NOR2X1 U1401 ( .A(BUSA[11]), .B(n1823), .Y(n1739) );
  NOR2X1 U1402 ( .A(n1707), .B(n1706), .Y(n1709) );
  NOR2X1 U1403 ( .A(n1800), .B(n1705), .Y(n1706) );
  NOR2X1 U1404 ( .A(BUSA[9]), .B(n1823), .Y(n1705) );
  NOR2X1 U1405 ( .A(n1779), .B(n1778), .Y(n1782) );
  NOR2X1 U1406 ( .A(n1800), .B(n1777), .Y(n1778) );
  NOR2X1 U1407 ( .A(BUSA[13]), .B(n1823), .Y(n1777) );
  OAI21XL U1408 ( .A0(n1441), .A1(n857), .B0(n1440), .Y(n1446) );
  OAI21XL U1409 ( .A0(n1474), .A1(n1163), .B0(n1443), .Y(n1445) );
  NOR2XL U1410 ( .A(n1350), .B(n873), .Y(n1364) );
  NOR2XL U1411 ( .A(n1346), .B(n874), .Y(n1366) );
  NOR2XL U1412 ( .A(n1350), .B(n874), .Y(n1241) );
  NOR2XL U1413 ( .A(n1422), .B(n874), .Y(n1257) );
  NOR2X1 U1414 ( .A(n1420), .B(n1163), .Y(n1365) );
  NOR2X1 U1415 ( .A(n1420), .B(n857), .Y(n1258) );
  NAND2X1 U1416 ( .A(n1330), .B(n1463), .Y(n1335) );
  NOR2XL U1417 ( .A(n1441), .B(n873), .Y(n1304) );
  NOR2XL U1418 ( .A(n1474), .B(n874), .Y(n1502) );
  NOR2XL U1419 ( .A(n1522), .B(n873), .Y(n1180) );
  NOR2XL U1420 ( .A(n1521), .B(n874), .Y(n1181) );
  NOR2XL U1421 ( .A(n1323), .B(n873), .Y(n1192) );
  NAND2X1 U1422 ( .A(n1308), .B(n1307), .Y(n1381) );
  NOR2X1 U1423 ( .A(n1422), .B(n857), .Y(n1306) );
  NAND2X1 U1424 ( .A(n1457), .B(n1464), .Y(n1373) );
  NOR2XL U1425 ( .A(n1418), .B(n873), .Y(n1255) );
  NAND2X1 U1426 ( .A(n1260), .B(n1259), .Y(n1345) );
  NOR2X1 U1427 ( .A(n1256), .B(n1255), .Y(n1260) );
  NAND4X1 U1428 ( .A(n1252), .B(n1426), .C(n1251), .D(n1250), .Y(n1430) );
  NAND2X1 U1429 ( .A(n1421), .B(n1521), .Y(n1251) );
  NAND2X1 U1430 ( .A(n1423), .B(n1474), .Y(n1250) );
  NOR2X1 U1431 ( .A(n1395), .B(n1485), .Y(n1217) );
  NAND2X1 U1432 ( .A(n1423), .B(n1350), .Y(n1351) );
  NOR2X1 U1433 ( .A(n1474), .B(n857), .Y(n1189) );
  NAND2X1 U1434 ( .A(n1191), .B(n1190), .Y(n1466) );
  NAND2X1 U1435 ( .A(n1196), .B(n1195), .Y(n1316) );
  NOR2XL U1436 ( .A(n1520), .B(n869), .Y(n1465) );
  NOR2X1 U1437 ( .A(n1406), .B(n1287), .Y(n1275) );
  NOR2XL U1438 ( .A(n1422), .B(n869), .Y(n1397) );
  NOR2XL U1439 ( .A(n1474), .B(n869), .Y(n1449) );
  NOR2XL U1440 ( .A(n1441), .B(n869), .Y(n1429) );
  NOR2X1 U1441 ( .A(n1758), .B(n847), .Y(n1753) );
  NOR2XL U1442 ( .A(n1406), .B(n874), .Y(n1194) );
  NOR2XL U1443 ( .A(n1722), .B(n847), .Y(n1718) );
  NOR2XL U1444 ( .A(n1689), .B(n847), .Y(n1684) );
  NOR2X1 U1445 ( .A(n1521), .B(n898), .Y(n1481) );
  NOR2BX1 U1446 ( .AN(n1466), .B(n1362), .Y(n1201) );
  CLKBUFX3 U1447 ( .A(n1143), .Y(n1139) );
  CLKBUFX3 U1448 ( .A(n1144), .Y(n1140) );
  CLKINVX1 U1449 ( .A(n1496), .Y(n1499) );
  AND2XL U1450 ( .A(n1482), .B(n874), .Y(n1279) );
  CLKBUFX3 U1451 ( .A(n1151), .Y(n1147) );
  CLKINVX1 U1452 ( .A(n1485), .Y(n1457) );
  NOR2X1 U1453 ( .A(n1406), .B(n1208), .Y(n1229) );
  AND2X2 U1454 ( .A(n1539), .B(n1851), .Y(n899) );
  CLKINVX1 U1455 ( .A(n899), .Y(n1856) );
  NOR2XL U1456 ( .A(n1346), .B(n873), .Y(n1239) );
  NAND2BX1 U1457 ( .AN(BUSA[0]), .B(n1174), .Y(n1565) );
  CLKINVX1 U1458 ( .A(n1464), .Y(n1292) );
  NAND2X1 U1459 ( .A(n1538), .B(n1543), .Y(n1547) );
  CLKBUFX3 U1460 ( .A(n1144), .Y(n1141) );
  CLKBUFX3 U1461 ( .A(n1144), .Y(n1142) );
  CLKBUFX3 U1462 ( .A(n1152), .Y(n1149) );
  CLKBUFX3 U1463 ( .A(n1152), .Y(n1148) );
  AOI21X1 U1464 ( .A0(N67), .A1(n1868), .B0(n1832), .Y(n1833) );
  NOR2X1 U1465 ( .A(n1831), .B(n1830), .Y(n1832) );
  AND3X2 U1466 ( .A(n918), .B(n1551), .C(n1550), .Y(n900) );
  INVX1 U1467 ( .A(n847), .Y(n1800) );
  CLKINVX1 U1468 ( .A(n1795), .Y(n1813) );
  AND2X2 U1469 ( .A(n919), .B(n1550), .Y(n901) );
  CLKINVX1 U1470 ( .A(n1757), .Y(n1820) );
  CLKINVX1 U1471 ( .A(n1814), .Y(n1860) );
  CLKINVX1 U1472 ( .A(BUSA[15]), .Y(n1861) );
  CLKBUFX3 U1473 ( .A(n1152), .Y(n1150) );
  AOI21X1 U1474 ( .A0(N73), .A1(n1868), .B0(n1715), .Y(n1716) );
  CLKINVX1 U1475 ( .A(n1835), .Y(n1717) );
  CLKINVX1 U1476 ( .A(n1837), .Y(n1752) );
  CLKINVX1 U1477 ( .A(n1839), .Y(n1789) );
  NOR2X1 U1478 ( .A(n1831), .B(n1732), .Y(n1733) );
  NOR2X1 U1479 ( .A(n1831), .B(n1770), .Y(n1771) );
  NOR2X1 U1480 ( .A(n1831), .B(n1808), .Y(n1809) );
  NOR2X1 U1481 ( .A(n1867), .B(n1866), .Y(n112) );
  CLKINVX1 U1482 ( .A(n129), .Y(n1831) );
  AND2X2 U1483 ( .A(n94), .B(n86), .Y(n902) );
  CLKINVX1 U1484 ( .A(n902), .Y(n121) );
  AND2X2 U1485 ( .A(n97), .B(n86), .Y(n903) );
  CLKINVX1 U1486 ( .A(n903), .Y(n123) );
  AND2X2 U1487 ( .A(n97), .B(n93), .Y(n904) );
  CLKINVX1 U1488 ( .A(n904), .Y(n95) );
  AND2X2 U1489 ( .A(n112), .B(n94), .Y(n905) );
  CLKINVX1 U1490 ( .A(n905), .Y(n110) );
  AND2X2 U1491 ( .A(n112), .B(n97), .Y(n906) );
  CLKINVX1 U1492 ( .A(n906), .Y(n113) );
  AND2X2 U1493 ( .A(n93), .B(n94), .Y(n907) );
  CLKINVX1 U1494 ( .A(n907), .Y(n91) );
  AND2X2 U1495 ( .A(n105), .B(n94), .Y(n908) );
  CLKINVX1 U1496 ( .A(n908), .Y(n103) );
  AND2X2 U1497 ( .A(n105), .B(n97), .Y(n909) );
  CLKINVX1 U1498 ( .A(n909), .Y(n106) );
  AND2X2 U1499 ( .A(n112), .B(n87), .Y(n910) );
  CLKINVX1 U1500 ( .A(n910), .Y(n115) );
  AND2X2 U1501 ( .A(n112), .B(n90), .Y(n911) );
  CLKINVX1 U1502 ( .A(n911), .Y(n118) );
  AND2X2 U1503 ( .A(n86), .B(n87), .Y(n912) );
  CLKINVX1 U1504 ( .A(n912), .Y(n69) );
  AND2X2 U1505 ( .A(n90), .B(n86), .Y(n913) );
  CLKINVX1 U1506 ( .A(n913), .Y(n88) );
  AND2X2 U1507 ( .A(n93), .B(n87), .Y(n914) );
  CLKINVX1 U1508 ( .A(n914), .Y(n98) );
  AND2X2 U1509 ( .A(n93), .B(n90), .Y(n915) );
  CLKINVX1 U1510 ( .A(n915), .Y(n100) );
  AND2X2 U1511 ( .A(n105), .B(n87), .Y(n916) );
  CLKINVX1 U1512 ( .A(n916), .Y(n108) );
  AND2X2 U1513 ( .A(n105), .B(n90), .Y(n917) );
  CLKINVX1 U1514 ( .A(n917), .Y(n126) );
  CLKINVX1 U1515 ( .A(n128), .Y(n1834) );
  CLKBUFX3 U1516 ( .A(n1000), .Y(n997) );
  CLKBUFX3 U1517 ( .A(n1000), .Y(n998) );
  CLKBUFX3 U1518 ( .A(n999), .Y(n994) );
  CLKBUFX3 U1519 ( .A(n999), .Y(n995) );
  CLKBUFX3 U1520 ( .A(n1000), .Y(n996) );
  CLKBUFX3 U1521 ( .A(n999), .Y(n993) );
  MXI4X1 U1522 ( .A(R12[1]), .B(R13[1]), .C(R14[1]), .D(R15[1]), .S0(n1138), 
        .S1(n1146), .Y(n1080) );
  MXI4X1 U1523 ( .A(R4[1]), .B(R5[1]), .C(R6[1]), .D(R7[1]), .S0(n1138), .S1(
        n1146), .Y(n1079) );
  MXI4X1 U1524 ( .A(R0[1]), .B(R1[1]), .C(R2[1]), .D(R3[1]), .S0(n1138), .S1(
        n1146), .Y(n1077) );
  MXI4X1 U1525 ( .A(R4[2]), .B(R5[2]), .C(R6[2]), .D(R7[2]), .S0(n1138), .S1(
        n1146), .Y(n1083) );
  MXI4X1 U1526 ( .A(R12[2]), .B(R13[2]), .C(R14[2]), .D(R15[2]), .S0(n1138), 
        .S1(n1146), .Y(n1084) );
  MXI4X1 U1527 ( .A(R0[2]), .B(R1[2]), .C(R2[2]), .D(R3[2]), .S0(n1138), .S1(
        n1146), .Y(n1081) );
  MXI4X1 U1528 ( .A(R4[3]), .B(R5[3]), .C(R6[3]), .D(R7[3]), .S0(n1138), .S1(
        n1146), .Y(n1087) );
  MXI4X1 U1529 ( .A(R12[3]), .B(R13[3]), .C(R14[3]), .D(R15[3]), .S0(n1138), 
        .S1(n1146), .Y(n1088) );
  MXI4X1 U1530 ( .A(R0[3]), .B(R1[3]), .C(R2[3]), .D(R3[3]), .S0(n1138), .S1(
        n1146), .Y(n1085) );
  MXI4X1 U1531 ( .A(R12[0]), .B(R13[0]), .C(R14[0]), .D(R15[0]), .S0(N57), 
        .S1(n1065), .Y(n1004) );
  MXI4X1 U1532 ( .A(R4[0]), .B(R5[0]), .C(R6[0]), .D(R7[0]), .S0(N57), .S1(
        n1065), .Y(n1003) );
  MXI2X4 U1533 ( .A(N109), .B(constant[6]), .S0(control[13]), .Y(n1441) );
  MXI4X2 U1534 ( .A(n1025), .B(n1026), .C(n1027), .D(n1028), .S0(N60), .S1(N59), .Y(N109) );
  MXI4X1 U1535 ( .A(R12[6]), .B(R13[6]), .C(R14[6]), .D(R15[6]), .S0(N57), 
        .S1(n1067), .Y(n1028) );
  MXI4X1 U1536 ( .A(R4[6]), .B(R5[6]), .C(R6[6]), .D(R7[6]), .S0(N57), .S1(
        n1067), .Y(n1027) );
  MXI4X2 U1537 ( .A(n1049), .B(n1050), .C(n1051), .D(n1052), .S0(N60), .S1(N59), .Y(N103) );
  NAND3X1 U1538 ( .A(n1202), .B(control[7]), .C(n1185), .Y(n1203) );
  MXI4X1 U1539 ( .A(R12[13]), .B(R13[13]), .C(R14[13]), .D(R15[13]), .S0(N57), 
        .S1(n1070), .Y(n1056) );
  MXI4X1 U1540 ( .A(R4[13]), .B(R5[13]), .C(R6[13]), .D(R7[13]), .S0(N57), 
        .S1(n1070), .Y(n1055) );
  NAND2X1 U1541 ( .A(n1415), .B(control[4]), .Y(n1455) );
  MXI4X1 U1542 ( .A(R4[15]), .B(R5[15]), .C(R6[15]), .D(R7[15]), .S0(N57), 
        .S1(n1070), .Y(n1063) );
  CLKBUFX3 U1543 ( .A(n1878), .Y(BUSA[0]) );
  MXI4X1 U1544 ( .A(n1073), .B(n1074), .C(n1075), .D(n1076), .S0(N64), .S1(N63), .Y(n1878) );
  MXI4X1 U1545 ( .A(R12[0]), .B(R13[0]), .C(R14[0]), .D(R15[0]), .S0(n1137), 
        .S1(n1145), .Y(n1076) );
  MXI4X1 U1546 ( .A(R4[0]), .B(R5[0]), .C(R6[0]), .D(R7[0]), .S0(n1137), .S1(
        n1145), .Y(n1075) );
  OR2X1 U1547 ( .A(n1406), .B(n1263), .Y(n1372) );
  NAND2X1 U1548 ( .A(n1264), .B(control[5]), .Y(n1263) );
  MXI4X1 U1549 ( .A(R0[0]), .B(R1[0]), .C(R2[0]), .D(R3[0]), .S0(N57), .S1(
        n1065), .Y(n1001) );
  MXI4X1 U1550 ( .A(R0[0]), .B(R1[0]), .C(R2[0]), .D(R3[0]), .S0(n1137), .S1(
        n1145), .Y(n1073) );
  MXI4X1 U1551 ( .A(R0[7]), .B(R1[7]), .C(R2[7]), .D(R3[7]), .S0(N57), .S1(
        n1068), .Y(n1029) );
  MXI4X1 U1552 ( .A(R0[10]), .B(R1[10]), .C(R2[10]), .D(R3[10]), .S0(N57), 
        .S1(n1069), .Y(n1041) );
  MXI4X1 U1553 ( .A(R0[11]), .B(R1[11]), .C(R2[11]), .D(R3[11]), .S0(N57), 
        .S1(n1069), .Y(n1045) );
  MXI4X1 U1554 ( .A(R8[0]), .B(R9[0]), .C(R10[0]), .D(R11[0]), .S0(N57), .S1(
        n1065), .Y(n1002) );
  MXI4X1 U1555 ( .A(R8[0]), .B(R9[0]), .C(R10[0]), .D(R11[0]), .S0(n1137), 
        .S1(n1145), .Y(n1074) );
  MXI4X1 U1556 ( .A(R8[7]), .B(R9[7]), .C(R10[7]), .D(R11[7]), .S0(N57), .S1(
        n1068), .Y(n1030) );
  MXI4X1 U1557 ( .A(R8[10]), .B(R9[10]), .C(R10[10]), .D(R11[10]), .S0(N57), 
        .S1(n1069), .Y(n1042) );
  MXI4X1 U1558 ( .A(R8[11]), .B(R9[11]), .C(R10[11]), .D(R11[11]), .S0(N57), 
        .S1(n1069), .Y(n1046) );
  MXI4X1 U1559 ( .A(R8[2]), .B(R9[2]), .C(R10[2]), .D(R11[2]), .S0(n1138), 
        .S1(n1146), .Y(n1082) );
  MXI4X1 U1560 ( .A(R8[3]), .B(R9[3]), .C(R10[3]), .D(R11[3]), .S0(n1138), 
        .S1(n1146), .Y(n1086) );
  CLKBUFX3 U1561 ( .A(N62), .Y(n1151) );
  MXI4X1 U1562 ( .A(R4[7]), .B(R5[7]), .C(R6[7]), .D(R7[7]), .S0(n1140), .S1(
        n1148), .Y(n1103) );
  MXI4X1 U1563 ( .A(R12[7]), .B(R13[7]), .C(R14[7]), .D(R15[7]), .S0(n1140), 
        .S1(n1148), .Y(n1104) );
  MXI4X1 U1564 ( .A(R0[7]), .B(R1[7]), .C(R2[7]), .D(R3[7]), .S0(n1140), .S1(
        n1148), .Y(n1101) );
  MXI4X1 U1565 ( .A(R4[4]), .B(R5[4]), .C(R6[4]), .D(R7[4]), .S0(n1139), .S1(
        n1147), .Y(n1091) );
  MXI4X1 U1566 ( .A(R12[4]), .B(R13[4]), .C(R14[4]), .D(R15[4]), .S0(n1139), 
        .S1(n1147), .Y(n1092) );
  MXI4X1 U1567 ( .A(R0[4]), .B(R1[4]), .C(R2[4]), .D(R3[4]), .S0(n1139), .S1(
        n1147), .Y(n1089) );
  MXI4X1 U1568 ( .A(R4[5]), .B(R5[5]), .C(R6[5]), .D(R7[5]), .S0(n1139), .S1(
        n1147), .Y(n1095) );
  MXI4X1 U1569 ( .A(R12[5]), .B(R13[5]), .C(R14[5]), .D(R15[5]), .S0(n1139), 
        .S1(n1147), .Y(n1096) );
  MXI4X1 U1570 ( .A(R0[5]), .B(R1[5]), .C(R2[5]), .D(R3[5]), .S0(n1139), .S1(
        n1147), .Y(n1093) );
  MXI4X1 U1571 ( .A(R4[6]), .B(R5[6]), .C(R6[6]), .D(R7[6]), .S0(n1139), .S1(
        n1147), .Y(n1099) );
  MXI4X1 U1572 ( .A(R12[6]), .B(R13[6]), .C(R14[6]), .D(R15[6]), .S0(n1139), 
        .S1(n1147), .Y(n1100) );
  MXI4X1 U1573 ( .A(R0[6]), .B(R1[6]), .C(R2[6]), .D(R3[6]), .S0(n1139), .S1(
        n1147), .Y(n1097) );
  OAI22XL U1574 ( .A0(control[4]), .A1(n1387), .B0(n1384), .B1(n1328), .Y(
        n1462) );
  NAND3BX1 U1575 ( .AN(control[8]), .B(n1221), .C(control[6]), .Y(n1222) );
  NAND4X1 U1576 ( .A(n1249), .B(n874), .C(n1248), .D(n1247), .Y(n1496) );
  NAND2X1 U1577 ( .A(control[4]), .B(n1463), .Y(n1362) );
  NAND2X1 U1578 ( .A(control[3]), .B(n1406), .Y(n1276) );
  CLKINVX1 U1579 ( .A(control[6]), .Y(n1185) );
  CLKINVX1 U1580 ( .A(control[7]), .Y(n1221) );
  MXI4X1 U1581 ( .A(R8[4]), .B(R9[4]), .C(R10[4]), .D(R11[4]), .S0(n1139), 
        .S1(n1147), .Y(n1090) );
  MXI4X1 U1582 ( .A(R8[5]), .B(R9[5]), .C(R10[5]), .D(R11[5]), .S0(n1139), 
        .S1(n1147), .Y(n1094) );
  MXI4X1 U1583 ( .A(R8[6]), .B(R9[6]), .C(R10[6]), .D(R11[6]), .S0(n1139), 
        .S1(n1147), .Y(n1098) );
  MXI4X1 U1584 ( .A(R8[7]), .B(R9[7]), .C(R10[7]), .D(R11[7]), .S0(n1140), 
        .S1(n1148), .Y(n1102) );
  CLKBUFX3 U1585 ( .A(N61), .Y(n1144) );
  CLKINVX1 U1586 ( .A(control[8]), .Y(n1183) );
  NAND3X1 U1587 ( .A(n918), .B(control[11]), .C(n1551), .Y(n1851) );
  NAND3X1 U1588 ( .A(n1544), .B(control[11]), .C(n1551), .Y(n1539) );
  CLKBUFX3 U1589 ( .A(n1875), .Y(BUSA[10]) );
  MXI4X1 U1590 ( .A(n1113), .B(n1114), .C(n1115), .D(n1116), .S0(N64), .S1(N63), .Y(n1875) );
  MXI4X1 U1591 ( .A(R4[10]), .B(R5[10]), .C(R6[10]), .D(R7[10]), .S0(n1141), 
        .S1(n1149), .Y(n1115) );
  MXI4X1 U1592 ( .A(R12[10]), .B(R13[10]), .C(R14[10]), .D(R15[10]), .S0(n1141), .S1(n1149), .Y(n1116) );
  CLKBUFX3 U1593 ( .A(n1873), .Y(BUSA[12]) );
  MXI4X1 U1594 ( .A(n1121), .B(n1122), .C(n1123), .D(n1124), .S0(N64), .S1(N63), .Y(n1873) );
  MXI4X1 U1595 ( .A(R4[12]), .B(R5[12]), .C(R6[12]), .D(R7[12]), .S0(n1141), 
        .S1(n1149), .Y(n1123) );
  MXI4X1 U1596 ( .A(R12[12]), .B(R13[12]), .C(R14[12]), .D(R15[12]), .S0(n1141), .S1(n1149), .Y(n1124) );
  CLKBUFX3 U1597 ( .A(n1874), .Y(BUSA[11]) );
  MXI4X1 U1598 ( .A(n1117), .B(n1118), .C(n1119), .D(n1120), .S0(N64), .S1(N63), .Y(n1874) );
  MXI4X1 U1599 ( .A(R4[11]), .B(R5[11]), .C(R6[11]), .D(R7[11]), .S0(n1141), 
        .S1(n1149), .Y(n1119) );
  MXI4X1 U1600 ( .A(R12[11]), .B(R13[11]), .C(R14[11]), .D(R15[11]), .S0(n1141), .S1(n1149), .Y(n1120) );
  CLKBUFX3 U1601 ( .A(n1872), .Y(BUSA[13]) );
  MXI4X1 U1602 ( .A(n1125), .B(n1126), .C(n1127), .D(n1128), .S0(N64), .S1(N63), .Y(n1872) );
  MXI4X1 U1603 ( .A(R4[13]), .B(R5[13]), .C(R6[13]), .D(R7[13]), .S0(n1142), 
        .S1(n1150), .Y(n1127) );
  MXI4X1 U1604 ( .A(R12[13]), .B(R13[13]), .C(R14[13]), .D(R15[13]), .S0(n1142), .S1(n1150), .Y(n1128) );
  CLKBUFX3 U1605 ( .A(n1871), .Y(BUSA[14]) );
  MXI4X1 U1606 ( .A(n1129), .B(n1130), .C(n1131), .D(n1132), .S0(N64), .S1(N63), .Y(n1871) );
  MXI4X1 U1607 ( .A(R4[14]), .B(R5[14]), .C(R6[14]), .D(R7[14]), .S0(n1142), 
        .S1(n1150), .Y(n1131) );
  MXI4X1 U1608 ( .A(R12[14]), .B(R13[14]), .C(R14[14]), .D(R15[14]), .S0(n1142), .S1(n1150), .Y(n1132) );
  CLKBUFX3 U1609 ( .A(n1877), .Y(BUSA[8]) );
  MXI4X1 U1610 ( .A(n1105), .B(n1106), .C(n1107), .D(n1108), .S0(N64), .S1(N63), .Y(n1877) );
  MXI4X1 U1611 ( .A(R4[8]), .B(R5[8]), .C(R6[8]), .D(R7[8]), .S0(n1140), .S1(
        n1148), .Y(n1107) );
  MXI4X1 U1612 ( .A(R12[8]), .B(R13[8]), .C(R14[8]), .D(R15[8]), .S0(n1140), 
        .S1(n1148), .Y(n1108) );
  CLKBUFX3 U1613 ( .A(n1876), .Y(BUSA[9]) );
  MXI4X1 U1614 ( .A(n1109), .B(n1110), .C(n1111), .D(n1112), .S0(N64), .S1(N63), .Y(n1876) );
  MXI4X1 U1615 ( .A(R4[9]), .B(R5[9]), .C(R6[9]), .D(R7[9]), .S0(n1140), .S1(
        n1148), .Y(n1111) );
  MXI4X1 U1616 ( .A(R12[9]), .B(R13[9]), .C(R14[9]), .D(R15[9]), .S0(n1140), 
        .S1(n1148), .Y(n1112) );
  CLKINVX1 U1617 ( .A(control[10]), .Y(n1551) );
  AND2X2 U1618 ( .A(control[9]), .B(n1538), .Y(n918) );
  MXI4X1 U1619 ( .A(R0[8]), .B(R1[8]), .C(R2[8]), .D(R3[8]), .S0(n1140), .S1(
        n1148), .Y(n1105) );
  MXI4X1 U1620 ( .A(R0[9]), .B(R1[9]), .C(R2[9]), .D(R3[9]), .S0(n1140), .S1(
        n1148), .Y(n1109) );
  MXI4X1 U1621 ( .A(R0[10]), .B(R1[10]), .C(R2[10]), .D(R3[10]), .S0(n1141), 
        .S1(n1149), .Y(n1113) );
  MXI4X1 U1622 ( .A(R0[11]), .B(R1[11]), .C(R2[11]), .D(R3[11]), .S0(n1141), 
        .S1(n1149), .Y(n1117) );
  MXI4X1 U1623 ( .A(R0[12]), .B(R1[12]), .C(R2[12]), .D(R3[12]), .S0(n1141), 
        .S1(n1149), .Y(n1121) );
  MXI4X1 U1624 ( .A(R0[13]), .B(R1[13]), .C(R2[13]), .D(R3[13]), .S0(n1142), 
        .S1(n1150), .Y(n1125) );
  MXI4X1 U1625 ( .A(R0[14]), .B(R1[14]), .C(R2[14]), .D(R3[14]), .S0(n1142), 
        .S1(n1150), .Y(n1129) );
  MXI4X1 U1626 ( .A(R8[8]), .B(R9[8]), .C(R10[8]), .D(R11[8]), .S0(n1140), 
        .S1(n1148), .Y(n1106) );
  MXI4X1 U1627 ( .A(R8[9]), .B(R9[9]), .C(R10[9]), .D(R11[9]), .S0(n1140), 
        .S1(n1148), .Y(n1110) );
  MXI4X1 U1628 ( .A(R8[10]), .B(R9[10]), .C(R10[10]), .D(R11[10]), .S0(n1141), 
        .S1(n1149), .Y(n1114) );
  MXI4X1 U1629 ( .A(R8[11]), .B(R9[11]), .C(R10[11]), .D(R11[11]), .S0(n1141), 
        .S1(n1149), .Y(n1118) );
  MXI4X1 U1630 ( .A(R8[12]), .B(R9[12]), .C(R10[12]), .D(R11[12]), .S0(n1141), 
        .S1(n1149), .Y(n1122) );
  MXI4X1 U1631 ( .A(R8[13]), .B(R9[13]), .C(R10[13]), .D(R11[13]), .S0(n1142), 
        .S1(n1150), .Y(n1126) );
  MXI4X1 U1632 ( .A(R8[14]), .B(R9[14]), .C(R10[14]), .D(R11[14]), .S0(n1142), 
        .S1(n1150), .Y(n1130) );
  CLKINVX1 U1633 ( .A(control[12]), .Y(n1538) );
  CLKBUFX3 U1634 ( .A(N62), .Y(n1152) );
  CLKINVX1 U1635 ( .A(control[9]), .Y(n1543) );
  AOI21X1 U1636 ( .A0(n1548), .A1(n1547), .B0(control[10]), .Y(n1549) );
  NAND2X1 U1637 ( .A(control[12]), .B(control[9]), .Y(n1548) );
  NAND3X1 U1638 ( .A(control[10]), .B(control[11]), .C(n1544), .Y(n1814) );
  NAND3X1 U1639 ( .A(n1544), .B(control[10]), .C(n1550), .Y(n1811) );
  OAI22XL U1640 ( .A0(n110), .A1(n837), .B0(n339), .B1(n905), .Y(n595) );
  OAI22XL U1641 ( .A0(n113), .A1(n837), .B0(n355), .B1(n906), .Y(n611) );
  OAI22XL U1642 ( .A0(n115), .A1(n837), .B0(n371), .B1(n910), .Y(n627) );
  OAI22XL U1643 ( .A0(n118), .A1(n837), .B0(n387), .B1(n911), .Y(n643) );
  OAI22XL U1644 ( .A0(n121), .A1(n837), .B0(n403), .B1(n902), .Y(n659) );
  OAI22XL U1645 ( .A0(n123), .A1(n837), .B0(n419), .B1(n903), .Y(n675) );
  OAI22XL U1646 ( .A0(n69), .A1(n837), .B0(n435), .B1(n912), .Y(n691) );
  OAI22XL U1647 ( .A0(n88), .A1(n837), .B0(n451), .B1(n913), .Y(n707) );
  OAI22XL U1648 ( .A0(n91), .A1(n837), .B0(n467), .B1(n907), .Y(n723) );
  OAI22XL U1649 ( .A0(n95), .A1(n837), .B0(n483), .B1(n904), .Y(n739) );
  OAI22XL U1650 ( .A0(n98), .A1(n837), .B0(n499), .B1(n914), .Y(n755) );
  OAI22XL U1651 ( .A0(n100), .A1(n837), .B0(n515), .B1(n915), .Y(n771) );
  OAI22XL U1652 ( .A0(n103), .A1(n837), .B0(n531), .B1(n908), .Y(n787) );
  OAI22XL U1653 ( .A0(n106), .A1(n837), .B0(n547), .B1(n909), .Y(n803) );
  OAI22XL U1654 ( .A0(n108), .A1(n837), .B0(n563), .B1(n916), .Y(n819) );
  OAI22XL U1655 ( .A0(n126), .A1(n837), .B0(n579), .B1(n917), .Y(n835) );
  CLKINVX1 U1656 ( .A(n1542), .Y(n1545) );
  NAND3BX1 U1657 ( .AN(control[11]), .B(control[10]), .C(control[12]), .Y(
        n1542) );
  CLKBUFX3 U1658 ( .A(n1870), .Y(BUSA[15]) );
  MXI4X1 U1659 ( .A(n1133), .B(n1134), .C(n1135), .D(n1136), .S0(N64), .S1(N63), .Y(n1870) );
  MXI4X1 U1660 ( .A(R12[15]), .B(R13[15]), .C(R14[15]), .D(R15[15]), .S0(n1142), .S1(n1150), .Y(n1136) );
  MXI4X1 U1661 ( .A(R4[15]), .B(R5[15]), .C(R6[15]), .D(R7[15]), .S0(n1142), 
        .S1(n1150), .Y(n1135) );
  AND2X2 U1662 ( .A(n918), .B(control[10]), .Y(n919) );
  CLKINVX1 U1663 ( .A(control[11]), .Y(n1550) );
  XOR2X1 U1664 ( .A(control[9]), .B(control[11]), .Y(n920) );
  MXI4X1 U1665 ( .A(R0[15]), .B(R1[15]), .C(R2[15]), .D(R3[15]), .S0(n1142), 
        .S1(n1150), .Y(n1133) );
  MXI4X1 U1666 ( .A(R8[15]), .B(R9[15]), .C(R10[15]), .D(R11[15]), .S0(n1142), 
        .S1(n1150), .Y(n1134) );
  OAI22XL U1667 ( .A0(n1170), .A1(n110), .B0(n330), .B1(n905), .Y(n586) );
  OAI22XL U1668 ( .A0(n1171), .A1(n110), .B0(n331), .B1(n905), .Y(n587) );
  OAI22XL U1669 ( .A0(n1172), .A1(n110), .B0(n332), .B1(n905), .Y(n588) );
  OAI22XL U1670 ( .A0(n110), .A1(n838), .B0(n333), .B1(n905), .Y(n589) );
  OAI22XL U1671 ( .A0(n110), .A1(n864), .B0(n334), .B1(n905), .Y(n590) );
  OAI22XL U1672 ( .A0(n110), .A1(n860), .B0(n335), .B1(n905), .Y(n591) );
  OAI22XL U1673 ( .A0(n110), .A1(n866), .B0(n336), .B1(n905), .Y(n592) );
  OAI22XL U1674 ( .A0(n110), .A1(n862), .B0(n337), .B1(n905), .Y(n593) );
  OAI22XL U1675 ( .A0(n110), .A1(n858), .B0(n338), .B1(n905), .Y(n594) );
  OAI22XL U1676 ( .A0(n1170), .A1(n113), .B0(n346), .B1(n906), .Y(n602) );
  OAI22XL U1677 ( .A0(n1171), .A1(n113), .B0(n347), .B1(n906), .Y(n603) );
  OAI22XL U1678 ( .A0(n1172), .A1(n113), .B0(n348), .B1(n906), .Y(n604) );
  OAI22XL U1679 ( .A0(n113), .A1(n838), .B0(n349), .B1(n906), .Y(n605) );
  OAI22XL U1680 ( .A0(n113), .A1(n864), .B0(n350), .B1(n906), .Y(n606) );
  OAI22XL U1681 ( .A0(n113), .A1(n860), .B0(n351), .B1(n906), .Y(n607) );
  OAI22XL U1682 ( .A0(n113), .A1(n866), .B0(n352), .B1(n906), .Y(n608) );
  OAI22XL U1683 ( .A0(n113), .A1(n862), .B0(n353), .B1(n906), .Y(n609) );
  OAI22XL U1684 ( .A0(n113), .A1(n858), .B0(n354), .B1(n906), .Y(n610) );
  OAI22XL U1685 ( .A0(n1170), .A1(n115), .B0(n362), .B1(n910), .Y(n618) );
  OAI22XL U1686 ( .A0(n1171), .A1(n115), .B0(n363), .B1(n910), .Y(n619) );
  OAI22XL U1687 ( .A0(n1172), .A1(n115), .B0(n364), .B1(n910), .Y(n620) );
  OAI22XL U1688 ( .A0(n115), .A1(n838), .B0(n365), .B1(n910), .Y(n621) );
  OAI22XL U1689 ( .A0(n115), .A1(n864), .B0(n366), .B1(n910), .Y(n622) );
  OAI22XL U1690 ( .A0(n115), .A1(n860), .B0(n367), .B1(n910), .Y(n623) );
  OAI22XL U1691 ( .A0(n115), .A1(n866), .B0(n368), .B1(n910), .Y(n624) );
  OAI22XL U1692 ( .A0(n115), .A1(n862), .B0(n369), .B1(n910), .Y(n625) );
  OAI22XL U1693 ( .A0(n115), .A1(n858), .B0(n370), .B1(n910), .Y(n626) );
  OAI22XL U1694 ( .A0(n1170), .A1(n118), .B0(n378), .B1(n911), .Y(n634) );
  OAI22XL U1695 ( .A0(n1171), .A1(n118), .B0(n379), .B1(n911), .Y(n635) );
  OAI22XL U1696 ( .A0(n1172), .A1(n118), .B0(n380), .B1(n911), .Y(n636) );
  OAI22XL U1697 ( .A0(n118), .A1(n838), .B0(n381), .B1(n911), .Y(n637) );
  OAI22XL U1698 ( .A0(n118), .A1(n864), .B0(n382), .B1(n911), .Y(n638) );
  OAI22XL U1699 ( .A0(n118), .A1(n860), .B0(n383), .B1(n911), .Y(n639) );
  OAI22XL U1700 ( .A0(n118), .A1(n866), .B0(n384), .B1(n911), .Y(n640) );
  OAI22XL U1701 ( .A0(n118), .A1(n862), .B0(n385), .B1(n911), .Y(n641) );
  OAI22XL U1702 ( .A0(n118), .A1(n858), .B0(n386), .B1(n911), .Y(n642) );
  OAI22XL U1703 ( .A0(n1170), .A1(n121), .B0(n394), .B1(n902), .Y(n650) );
  OAI22XL U1704 ( .A0(n1171), .A1(n121), .B0(n395), .B1(n902), .Y(n651) );
  OAI22XL U1705 ( .A0(n1172), .A1(n121), .B0(n396), .B1(n902), .Y(n652) );
  OAI22XL U1706 ( .A0(n121), .A1(n838), .B0(n397), .B1(n902), .Y(n653) );
  OAI22XL U1707 ( .A0(n121), .A1(n864), .B0(n398), .B1(n902), .Y(n654) );
  OAI22XL U1708 ( .A0(n121), .A1(n860), .B0(n399), .B1(n902), .Y(n655) );
  OAI22XL U1709 ( .A0(n121), .A1(n866), .B0(n400), .B1(n902), .Y(n656) );
  OAI22XL U1710 ( .A0(n121), .A1(n862), .B0(n401), .B1(n902), .Y(n657) );
  OAI22XL U1711 ( .A0(n121), .A1(n858), .B0(n402), .B1(n902), .Y(n658) );
  OAI22XL U1712 ( .A0(n1170), .A1(n123), .B0(n410), .B1(n903), .Y(n666) );
  OAI22XL U1713 ( .A0(n1171), .A1(n123), .B0(n411), .B1(n903), .Y(n667) );
  OAI22XL U1714 ( .A0(n1172), .A1(n123), .B0(n412), .B1(n903), .Y(n668) );
  OAI22XL U1715 ( .A0(n123), .A1(n838), .B0(n413), .B1(n903), .Y(n669) );
  OAI22XL U1716 ( .A0(n123), .A1(n864), .B0(n414), .B1(n903), .Y(n670) );
  OAI22XL U1717 ( .A0(n123), .A1(n860), .B0(n415), .B1(n903), .Y(n671) );
  OAI22XL U1718 ( .A0(n123), .A1(n866), .B0(n416), .B1(n903), .Y(n672) );
  OAI22XL U1719 ( .A0(n123), .A1(n862), .B0(n417), .B1(n903), .Y(n673) );
  OAI22XL U1720 ( .A0(n123), .A1(n858), .B0(n418), .B1(n903), .Y(n674) );
  OAI22XL U1721 ( .A0(n1170), .A1(n69), .B0(n426), .B1(n912), .Y(n682) );
  OAI22XL U1722 ( .A0(n1171), .A1(n69), .B0(n427), .B1(n912), .Y(n683) );
  OAI22XL U1723 ( .A0(n1172), .A1(n69), .B0(n428), .B1(n912), .Y(n684) );
  OAI22XL U1724 ( .A0(n69), .A1(n838), .B0(n429), .B1(n912), .Y(n685) );
  OAI22XL U1725 ( .A0(n69), .A1(n864), .B0(n430), .B1(n912), .Y(n686) );
  OAI22XL U1726 ( .A0(n69), .A1(n860), .B0(n431), .B1(n912), .Y(n687) );
  OAI22XL U1727 ( .A0(n69), .A1(n866), .B0(n432), .B1(n912), .Y(n688) );
  OAI22XL U1728 ( .A0(n69), .A1(n862), .B0(n433), .B1(n912), .Y(n689) );
  OAI22XL U1729 ( .A0(n69), .A1(n858), .B0(n434), .B1(n912), .Y(n690) );
  OAI22XL U1730 ( .A0(n1170), .A1(n88), .B0(n442), .B1(n913), .Y(n698) );
  OAI22XL U1731 ( .A0(n1171), .A1(n88), .B0(n443), .B1(n913), .Y(n699) );
  OAI22XL U1732 ( .A0(n1172), .A1(n88), .B0(n444), .B1(n913), .Y(n700) );
  OAI22XL U1733 ( .A0(n88), .A1(n838), .B0(n445), .B1(n913), .Y(n701) );
  OAI22XL U1734 ( .A0(n88), .A1(n864), .B0(n446), .B1(n913), .Y(n702) );
  OAI22XL U1735 ( .A0(n88), .A1(n860), .B0(n447), .B1(n913), .Y(n703) );
  OAI22XL U1736 ( .A0(n88), .A1(n866), .B0(n448), .B1(n913), .Y(n704) );
  OAI22XL U1737 ( .A0(n88), .A1(n862), .B0(n449), .B1(n913), .Y(n705) );
  OAI22XL U1738 ( .A0(n88), .A1(n858), .B0(n450), .B1(n913), .Y(n706) );
  OAI22XL U1739 ( .A0(n1170), .A1(n91), .B0(n458), .B1(n907), .Y(n714) );
  OAI22XL U1740 ( .A0(n1171), .A1(n91), .B0(n459), .B1(n907), .Y(n715) );
  OAI22XL U1741 ( .A0(n1172), .A1(n91), .B0(n460), .B1(n907), .Y(n716) );
  OAI22XL U1742 ( .A0(n91), .A1(n838), .B0(n461), .B1(n907), .Y(n717) );
  OAI22XL U1743 ( .A0(n91), .A1(n864), .B0(n462), .B1(n907), .Y(n718) );
  OAI22XL U1744 ( .A0(n91), .A1(n860), .B0(n463), .B1(n907), .Y(n719) );
  OAI22XL U1745 ( .A0(n91), .A1(n866), .B0(n464), .B1(n907), .Y(n720) );
  OAI22XL U1746 ( .A0(n91), .A1(n862), .B0(n465), .B1(n907), .Y(n721) );
  OAI22XL U1747 ( .A0(n91), .A1(n858), .B0(n466), .B1(n907), .Y(n722) );
  OAI22XL U1748 ( .A0(n1170), .A1(n95), .B0(n474), .B1(n904), .Y(n730) );
  OAI22XL U1749 ( .A0(n1171), .A1(n95), .B0(n475), .B1(n904), .Y(n731) );
  OAI22XL U1750 ( .A0(n1172), .A1(n95), .B0(n476), .B1(n904), .Y(n732) );
  OAI22XL U1751 ( .A0(n95), .A1(n838), .B0(n477), .B1(n904), .Y(n733) );
  OAI22XL U1752 ( .A0(n95), .A1(n864), .B0(n478), .B1(n904), .Y(n734) );
  OAI22XL U1753 ( .A0(n95), .A1(n860), .B0(n479), .B1(n904), .Y(n735) );
  OAI22XL U1754 ( .A0(n95), .A1(n866), .B0(n480), .B1(n904), .Y(n736) );
  OAI22XL U1755 ( .A0(n95), .A1(n862), .B0(n481), .B1(n904), .Y(n737) );
  OAI22XL U1756 ( .A0(n95), .A1(n858), .B0(n482), .B1(n904), .Y(n738) );
  OAI22XL U1757 ( .A0(n1170), .A1(n98), .B0(n490), .B1(n914), .Y(n746) );
  OAI22XL U1758 ( .A0(n1171), .A1(n98), .B0(n491), .B1(n914), .Y(n747) );
  OAI22XL U1759 ( .A0(n1172), .A1(n98), .B0(n492), .B1(n914), .Y(n748) );
  OAI22XL U1760 ( .A0(n98), .A1(n838), .B0(n493), .B1(n914), .Y(n749) );
  OAI22XL U1761 ( .A0(n98), .A1(n864), .B0(n494), .B1(n914), .Y(n750) );
  OAI22XL U1762 ( .A0(n98), .A1(n860), .B0(n495), .B1(n914), .Y(n751) );
  OAI22XL U1763 ( .A0(n98), .A1(n866), .B0(n496), .B1(n914), .Y(n752) );
  OAI22XL U1764 ( .A0(n98), .A1(n862), .B0(n497), .B1(n914), .Y(n753) );
  OAI22XL U1765 ( .A0(n98), .A1(n858), .B0(n498), .B1(n914), .Y(n754) );
  OAI22XL U1766 ( .A0(n1170), .A1(n100), .B0(n506), .B1(n915), .Y(n762) );
  OAI22XL U1767 ( .A0(n1171), .A1(n100), .B0(n507), .B1(n915), .Y(n763) );
  OAI22XL U1768 ( .A0(n1172), .A1(n100), .B0(n508), .B1(n915), .Y(n764) );
  OAI22XL U1769 ( .A0(n100), .A1(n838), .B0(n509), .B1(n915), .Y(n765) );
  OAI22XL U1770 ( .A0(n100), .A1(n864), .B0(n510), .B1(n915), .Y(n766) );
  OAI22XL U1771 ( .A0(n100), .A1(n860), .B0(n511), .B1(n915), .Y(n767) );
  OAI22XL U1772 ( .A0(n100), .A1(n866), .B0(n512), .B1(n915), .Y(n768) );
  OAI22XL U1773 ( .A0(n100), .A1(n862), .B0(n513), .B1(n915), .Y(n769) );
  OAI22XL U1774 ( .A0(n100), .A1(n858), .B0(n514), .B1(n915), .Y(n770) );
  OAI22XL U1775 ( .A0(n1170), .A1(n103), .B0(n522), .B1(n908), .Y(n778) );
  OAI22XL U1776 ( .A0(n1171), .A1(n103), .B0(n523), .B1(n908), .Y(n779) );
  OAI22XL U1777 ( .A0(n1172), .A1(n103), .B0(n524), .B1(n908), .Y(n780) );
  OAI22XL U1778 ( .A0(n103), .A1(n838), .B0(n525), .B1(n908), .Y(n781) );
  OAI22XL U1779 ( .A0(n103), .A1(n864), .B0(n526), .B1(n908), .Y(n782) );
  OAI22XL U1780 ( .A0(n103), .A1(n860), .B0(n527), .B1(n908), .Y(n783) );
  OAI22XL U1781 ( .A0(n103), .A1(n866), .B0(n528), .B1(n908), .Y(n784) );
  OAI22XL U1782 ( .A0(n103), .A1(n862), .B0(n529), .B1(n908), .Y(n785) );
  OAI22XL U1783 ( .A0(n103), .A1(n858), .B0(n530), .B1(n908), .Y(n786) );
  OAI22XL U1784 ( .A0(n1170), .A1(n106), .B0(n538), .B1(n909), .Y(n794) );
  OAI22XL U1785 ( .A0(n1171), .A1(n106), .B0(n539), .B1(n909), .Y(n795) );
  OAI22XL U1786 ( .A0(n1172), .A1(n106), .B0(n540), .B1(n909), .Y(n796) );
  OAI22XL U1787 ( .A0(n106), .A1(n838), .B0(n541), .B1(n909), .Y(n797) );
  OAI22XL U1788 ( .A0(n106), .A1(n864), .B0(n542), .B1(n909), .Y(n798) );
  OAI22XL U1789 ( .A0(n106), .A1(n860), .B0(n543), .B1(n909), .Y(n799) );
  OAI22XL U1790 ( .A0(n106), .A1(n866), .B0(n544), .B1(n909), .Y(n800) );
  OAI22XL U1791 ( .A0(n106), .A1(n862), .B0(n545), .B1(n909), .Y(n801) );
  OAI22XL U1792 ( .A0(n106), .A1(n858), .B0(n546), .B1(n909), .Y(n802) );
  OAI22XL U1793 ( .A0(n1170), .A1(n108), .B0(n554), .B1(n916), .Y(n810) );
  OAI22XL U1794 ( .A0(n1171), .A1(n108), .B0(n555), .B1(n916), .Y(n811) );
  OAI22XL U1795 ( .A0(n1172), .A1(n108), .B0(n556), .B1(n916), .Y(n812) );
  OAI22XL U1796 ( .A0(n108), .A1(n838), .B0(n557), .B1(n916), .Y(n813) );
  OAI22XL U1797 ( .A0(n108), .A1(n864), .B0(n558), .B1(n916), .Y(n814) );
  OAI22XL U1798 ( .A0(n108), .A1(n860), .B0(n559), .B1(n916), .Y(n815) );
  OAI22XL U1799 ( .A0(n108), .A1(n866), .B0(n560), .B1(n916), .Y(n816) );
  OAI22XL U1800 ( .A0(n108), .A1(n862), .B0(n561), .B1(n916), .Y(n817) );
  OAI22XL U1801 ( .A0(n108), .A1(n858), .B0(n562), .B1(n916), .Y(n818) );
  OAI22XL U1802 ( .A0(n126), .A1(n838), .B0(n573), .B1(n917), .Y(n829) );
  OAI22XL U1803 ( .A0(n126), .A1(n864), .B0(n574), .B1(n917), .Y(n830) );
  OAI22XL U1804 ( .A0(n126), .A1(n860), .B0(n575), .B1(n917), .Y(n831) );
  OAI22XL U1805 ( .A0(n126), .A1(n866), .B0(n576), .B1(n917), .Y(n832) );
  OAI22XL U1806 ( .A0(n126), .A1(n862), .B0(n577), .B1(n917), .Y(n833) );
  OAI22XL U1807 ( .A0(n126), .A1(n858), .B0(n578), .B1(n917), .Y(n834) );
  OAI22XL U1808 ( .A0(n570), .A1(n917), .B0(n1170), .B1(n126), .Y(n826) );
  OAI22XL U1809 ( .A0(n571), .A1(n917), .B0(n1171), .B1(n126), .Y(n827) );
  OAI22XL U1810 ( .A0(n572), .A1(n917), .B0(n1172), .B1(n126), .Y(n828) );
  CLKBUFX3 U1811 ( .A(n73), .Y(n1170) );
  AOI222XL U1812 ( .A0(N76), .A1(n1868), .B0(n128), .B1(n52), .C0(data[6]), 
        .C1(n129), .Y(n73) );
  MXI4X1 U1813 ( .A(n945), .B(n946), .C(n947), .D(n948), .S0(N56), .S1(N55), 
        .Y(N76) );
  MXI4X1 U1814 ( .A(R12[6]), .B(R13[6]), .C(R14[6]), .D(R15[6]), .S0(n987), 
        .S1(n995), .Y(n948) );
  CLKBUFX3 U1815 ( .A(n72), .Y(n1171) );
  AOI222XL U1816 ( .A0(N75), .A1(n1868), .B0(n128), .B1(n53), .C0(data[7]), 
        .C1(n129), .Y(n72) );
  MXI4X1 U1817 ( .A(n949), .B(n950), .C(n951), .D(n952), .S0(N56), .S1(N55), 
        .Y(N75) );
  MXI4X1 U1818 ( .A(R12[7]), .B(R13[7]), .C(R14[7]), .D(R15[7]), .S0(n988), 
        .S1(n996), .Y(n952) );
  CLKBUFX3 U1819 ( .A(n71), .Y(n1172) );
  AOI222XL U1820 ( .A0(N74), .A1(n1868), .B0(n128), .B1(n54), .C0(data[8]), 
        .C1(n129), .Y(n71) );
  MXI4X1 U1821 ( .A(n953), .B(n954), .C(n955), .D(n956), .S0(N56), .S1(N55), 
        .Y(N74) );
  MXI4X1 U1822 ( .A(R12[8]), .B(R13[8]), .C(R14[8]), .D(R15[8]), .S0(n988), 
        .S1(n996), .Y(n956) );
  OAI22XL U1823 ( .A0(n1164), .A1(n110), .B0(n324), .B1(n905), .Y(n580) );
  OAI22XL U1824 ( .A0(n1165), .A1(n110), .B0(n325), .B1(n905), .Y(n581) );
  OAI22XL U1825 ( .A0(n1166), .A1(n110), .B0(n326), .B1(n905), .Y(n582) );
  OAI22XL U1826 ( .A0(n1167), .A1(n110), .B0(n327), .B1(n905), .Y(n583) );
  OAI22XL U1827 ( .A0(n1168), .A1(n110), .B0(n328), .B1(n905), .Y(n584) );
  OAI22XL U1828 ( .A0(n1169), .A1(n110), .B0(n329), .B1(n905), .Y(n585) );
  OAI22XL U1829 ( .A0(n1164), .A1(n113), .B0(n340), .B1(n906), .Y(n596) );
  OAI22XL U1830 ( .A0(n1165), .A1(n113), .B0(n341), .B1(n906), .Y(n597) );
  OAI22XL U1831 ( .A0(n1166), .A1(n113), .B0(n342), .B1(n906), .Y(n598) );
  OAI22XL U1832 ( .A0(n1167), .A1(n113), .B0(n343), .B1(n906), .Y(n599) );
  OAI22XL U1833 ( .A0(n1168), .A1(n113), .B0(n344), .B1(n906), .Y(n600) );
  OAI22XL U1834 ( .A0(n1169), .A1(n113), .B0(n345), .B1(n906), .Y(n601) );
  OAI22XL U1835 ( .A0(n1164), .A1(n115), .B0(n356), .B1(n910), .Y(n612) );
  OAI22XL U1836 ( .A0(n1165), .A1(n115), .B0(n357), .B1(n910), .Y(n613) );
  OAI22XL U1837 ( .A0(n1166), .A1(n115), .B0(n358), .B1(n910), .Y(n614) );
  OAI22XL U1838 ( .A0(n1167), .A1(n115), .B0(n359), .B1(n910), .Y(n615) );
  OAI22XL U1839 ( .A0(n1168), .A1(n115), .B0(n360), .B1(n910), .Y(n616) );
  OAI22XL U1840 ( .A0(n1169), .A1(n115), .B0(n361), .B1(n910), .Y(n617) );
  OAI22XL U1841 ( .A0(n1164), .A1(n118), .B0(n372), .B1(n911), .Y(n628) );
  OAI22XL U1842 ( .A0(n1165), .A1(n118), .B0(n373), .B1(n911), .Y(n629) );
  OAI22XL U1843 ( .A0(n1166), .A1(n118), .B0(n374), .B1(n911), .Y(n630) );
  OAI22XL U1844 ( .A0(n1167), .A1(n118), .B0(n375), .B1(n911), .Y(n631) );
  OAI22XL U1845 ( .A0(n1168), .A1(n118), .B0(n376), .B1(n911), .Y(n632) );
  OAI22XL U1846 ( .A0(n1169), .A1(n118), .B0(n377), .B1(n911), .Y(n633) );
  OAI22XL U1847 ( .A0(n1164), .A1(n121), .B0(n388), .B1(n902), .Y(n644) );
  OAI22XL U1848 ( .A0(n1165), .A1(n121), .B0(n389), .B1(n902), .Y(n645) );
  OAI22XL U1849 ( .A0(n1166), .A1(n121), .B0(n390), .B1(n902), .Y(n646) );
  OAI22XL U1850 ( .A0(n1167), .A1(n121), .B0(n391), .B1(n902), .Y(n647) );
  OAI22XL U1851 ( .A0(n1168), .A1(n121), .B0(n392), .B1(n902), .Y(n648) );
  OAI22XL U1852 ( .A0(n1169), .A1(n121), .B0(n393), .B1(n902), .Y(n649) );
  OAI22XL U1853 ( .A0(n1164), .A1(n123), .B0(n404), .B1(n903), .Y(n660) );
  OAI22XL U1854 ( .A0(n1165), .A1(n123), .B0(n405), .B1(n903), .Y(n661) );
  OAI22XL U1855 ( .A0(n1166), .A1(n123), .B0(n406), .B1(n903), .Y(n662) );
  OAI22XL U1856 ( .A0(n1167), .A1(n123), .B0(n407), .B1(n903), .Y(n663) );
  OAI22XL U1857 ( .A0(n1168), .A1(n123), .B0(n408), .B1(n903), .Y(n664) );
  OAI22XL U1858 ( .A0(n1169), .A1(n123), .B0(n409), .B1(n903), .Y(n665) );
  OAI22XL U1859 ( .A0(n1164), .A1(n69), .B0(n420), .B1(n912), .Y(n676) );
  OAI22XL U1860 ( .A0(n1165), .A1(n69), .B0(n421), .B1(n912), .Y(n677) );
  OAI22XL U1861 ( .A0(n1166), .A1(n69), .B0(n422), .B1(n912), .Y(n678) );
  OAI22XL U1862 ( .A0(n1167), .A1(n69), .B0(n423), .B1(n912), .Y(n679) );
  OAI22XL U1863 ( .A0(n1168), .A1(n69), .B0(n424), .B1(n912), .Y(n680) );
  OAI22XL U1864 ( .A0(n1169), .A1(n69), .B0(n425), .B1(n912), .Y(n681) );
  OAI22XL U1865 ( .A0(n1164), .A1(n88), .B0(n436), .B1(n913), .Y(n692) );
  OAI22XL U1866 ( .A0(n1165), .A1(n88), .B0(n437), .B1(n913), .Y(n693) );
  OAI22XL U1867 ( .A0(n1166), .A1(n88), .B0(n438), .B1(n913), .Y(n694) );
  OAI22XL U1868 ( .A0(n1167), .A1(n88), .B0(n439), .B1(n913), .Y(n695) );
  OAI22XL U1869 ( .A0(n1168), .A1(n88), .B0(n440), .B1(n913), .Y(n696) );
  OAI22XL U1870 ( .A0(n1169), .A1(n88), .B0(n441), .B1(n913), .Y(n697) );
  OAI22XL U1871 ( .A0(n1164), .A1(n91), .B0(n452), .B1(n907), .Y(n708) );
  OAI22XL U1872 ( .A0(n1165), .A1(n91), .B0(n453), .B1(n907), .Y(n709) );
  OAI22XL U1873 ( .A0(n1166), .A1(n91), .B0(n454), .B1(n907), .Y(n710) );
  OAI22XL U1874 ( .A0(n1167), .A1(n91), .B0(n455), .B1(n907), .Y(n711) );
  OAI22XL U1875 ( .A0(n1168), .A1(n91), .B0(n456), .B1(n907), .Y(n712) );
  OAI22XL U1876 ( .A0(n1169), .A1(n91), .B0(n457), .B1(n907), .Y(n713) );
  OAI22XL U1877 ( .A0(n1164), .A1(n95), .B0(n468), .B1(n904), .Y(n724) );
  OAI22XL U1878 ( .A0(n1165), .A1(n95), .B0(n469), .B1(n904), .Y(n725) );
  OAI22XL U1879 ( .A0(n1166), .A1(n95), .B0(n470), .B1(n904), .Y(n726) );
  OAI22XL U1880 ( .A0(n1167), .A1(n95), .B0(n471), .B1(n904), .Y(n727) );
  OAI22XL U1881 ( .A0(n1168), .A1(n95), .B0(n472), .B1(n904), .Y(n728) );
  OAI22XL U1882 ( .A0(n1169), .A1(n95), .B0(n473), .B1(n904), .Y(n729) );
  OAI22XL U1883 ( .A0(n1164), .A1(n98), .B0(n484), .B1(n914), .Y(n740) );
  OAI22XL U1884 ( .A0(n1165), .A1(n98), .B0(n485), .B1(n914), .Y(n741) );
  OAI22XL U1885 ( .A0(n1166), .A1(n98), .B0(n486), .B1(n914), .Y(n742) );
  OAI22XL U1886 ( .A0(n1167), .A1(n98), .B0(n487), .B1(n914), .Y(n743) );
  OAI22XL U1887 ( .A0(n1168), .A1(n98), .B0(n488), .B1(n914), .Y(n744) );
  OAI22XL U1888 ( .A0(n1169), .A1(n98), .B0(n489), .B1(n914), .Y(n745) );
  OAI22XL U1889 ( .A0(n1164), .A1(n100), .B0(n500), .B1(n915), .Y(n756) );
  OAI22XL U1890 ( .A0(n1165), .A1(n100), .B0(n501), .B1(n915), .Y(n757) );
  OAI22XL U1891 ( .A0(n1166), .A1(n100), .B0(n502), .B1(n915), .Y(n758) );
  OAI22XL U1892 ( .A0(n1167), .A1(n100), .B0(n503), .B1(n915), .Y(n759) );
  OAI22XL U1893 ( .A0(n1168), .A1(n100), .B0(n504), .B1(n915), .Y(n760) );
  OAI22XL U1894 ( .A0(n1169), .A1(n100), .B0(n505), .B1(n915), .Y(n761) );
  OAI22XL U1895 ( .A0(n1164), .A1(n103), .B0(n516), .B1(n908), .Y(n772) );
  OAI22XL U1896 ( .A0(n1165), .A1(n103), .B0(n517), .B1(n908), .Y(n773) );
  OAI22XL U1897 ( .A0(n1166), .A1(n103), .B0(n518), .B1(n908), .Y(n774) );
  OAI22XL U1898 ( .A0(n1167), .A1(n103), .B0(n519), .B1(n908), .Y(n775) );
  OAI22XL U1899 ( .A0(n1168), .A1(n103), .B0(n520), .B1(n908), .Y(n776) );
  OAI22XL U1900 ( .A0(n1169), .A1(n103), .B0(n521), .B1(n908), .Y(n777) );
  OAI22XL U1901 ( .A0(n1164), .A1(n106), .B0(n532), .B1(n909), .Y(n788) );
  OAI22XL U1902 ( .A0(n1165), .A1(n106), .B0(n533), .B1(n909), .Y(n789) );
  OAI22XL U1903 ( .A0(n1166), .A1(n106), .B0(n534), .B1(n909), .Y(n790) );
  OAI22XL U1904 ( .A0(n1167), .A1(n106), .B0(n535), .B1(n909), .Y(n791) );
  OAI22XL U1905 ( .A0(n1168), .A1(n106), .B0(n536), .B1(n909), .Y(n792) );
  OAI22XL U1906 ( .A0(n1169), .A1(n106), .B0(n537), .B1(n909), .Y(n793) );
  OAI22XL U1907 ( .A0(n1164), .A1(n108), .B0(n548), .B1(n916), .Y(n804) );
  OAI22XL U1908 ( .A0(n1165), .A1(n108), .B0(n549), .B1(n916), .Y(n805) );
  OAI22XL U1909 ( .A0(n1166), .A1(n108), .B0(n550), .B1(n916), .Y(n806) );
  OAI22XL U1910 ( .A0(n1167), .A1(n108), .B0(n551), .B1(n916), .Y(n807) );
  OAI22XL U1911 ( .A0(n1168), .A1(n108), .B0(n552), .B1(n916), .Y(n808) );
  OAI22XL U1912 ( .A0(n1169), .A1(n108), .B0(n553), .B1(n916), .Y(n809) );
  OAI22XL U1913 ( .A0(n564), .A1(n917), .B0(n1164), .B1(n126), .Y(n820) );
  OAI22XL U1914 ( .A0(n565), .A1(n917), .B0(n1165), .B1(n126), .Y(n821) );
  OAI22XL U1915 ( .A0(n566), .A1(n917), .B0(n1166), .B1(n126), .Y(n822) );
  OAI22XL U1916 ( .A0(n567), .A1(n917), .B0(n1167), .B1(n126), .Y(n823) );
  OAI22XL U1917 ( .A0(n568), .A1(n917), .B0(n1168), .B1(n126), .Y(n824) );
  OAI22XL U1918 ( .A0(n569), .A1(n917), .B0(n1169), .B1(n126), .Y(n825) );
  CLKBUFX3 U1919 ( .A(n85), .Y(n1164) );
  AOI222XL U1920 ( .A0(N82), .A1(n1868), .B0(n128), .B1(n41), .C0(data[0]), 
        .C1(n129), .Y(n85) );
  MXI4X1 U1921 ( .A(n921), .B(n922), .C(n923), .D(n924), .S0(N56), .S1(N55), 
        .Y(N82) );
  MXI4X1 U1922 ( .A(R12[0]), .B(R13[0]), .C(R14[0]), .D(R15[0]), .S0(n985), 
        .S1(n993), .Y(n924) );
  CLKBUFX3 U1923 ( .A(n78), .Y(n1165) );
  AOI222XL U1924 ( .A0(N81), .A1(n1868), .B0(n128), .B1(n47), .C0(data[1]), 
        .C1(n129), .Y(n78) );
  MXI4X1 U1925 ( .A(n925), .B(n926), .C(n927), .D(n928), .S0(N56), .S1(N55), 
        .Y(N81) );
  MXI4X1 U1926 ( .A(R12[1]), .B(R13[1]), .C(R14[1]), .D(R15[1]), .S0(n986), 
        .S1(n994), .Y(n928) );
  CLKBUFX3 U1927 ( .A(n77), .Y(n1166) );
  AOI222XL U1928 ( .A0(N80), .A1(n1868), .B0(n128), .B1(n48), .C0(data[2]), 
        .C1(n129), .Y(n77) );
  MXI4X1 U1929 ( .A(n929), .B(n930), .C(n931), .D(n932), .S0(N56), .S1(N55), 
        .Y(N80) );
  MXI4X1 U1930 ( .A(R12[2]), .B(R13[2]), .C(R14[2]), .D(R15[2]), .S0(n986), 
        .S1(n994), .Y(n932) );
  CLKBUFX3 U1931 ( .A(n76), .Y(n1167) );
  AOI222XL U1932 ( .A0(N79), .A1(n1868), .B0(n128), .B1(n49), .C0(data[3]), 
        .C1(n129), .Y(n76) );
  MXI4X1 U1933 ( .A(n933), .B(n934), .C(n935), .D(n936), .S0(N56), .S1(N55), 
        .Y(N79) );
  MXI4X1 U1934 ( .A(R12[3]), .B(R13[3]), .C(R14[3]), .D(R15[3]), .S0(n986), 
        .S1(n994), .Y(n936) );
  CLKBUFX3 U1935 ( .A(n75), .Y(n1168) );
  AOI222XL U1936 ( .A0(N78), .A1(n1868), .B0(n128), .B1(n50), .C0(data[4]), 
        .C1(n129), .Y(n75) );
  MXI4X1 U1937 ( .A(n937), .B(n938), .C(n939), .D(n940), .S0(N56), .S1(N55), 
        .Y(N78) );
  MXI4X1 U1938 ( .A(R12[4]), .B(R13[4]), .C(R14[4]), .D(R15[4]), .S0(n987), 
        .S1(n995), .Y(n940) );
  CLKBUFX3 U1939 ( .A(n74), .Y(n1169) );
  AOI222XL U1940 ( .A0(N77), .A1(n1868), .B0(n128), .B1(n51), .C0(data[5]), 
        .C1(n129), .Y(n74) );
  MXI4X1 U1941 ( .A(n941), .B(n942), .C(n943), .D(n944), .S0(N56), .S1(N55), 
        .Y(N77) );
  MXI4X1 U1942 ( .A(R12[5]), .B(R13[5]), .C(R14[5]), .D(R15[5]), .S0(n987), 
        .S1(n995), .Y(n944) );
  MXI4X1 U1943 ( .A(n957), .B(n958), .C(n959), .D(n960), .S0(N56), .S1(N55), 
        .Y(N73) );
  MXI4X1 U1944 ( .A(R12[9]), .B(R13[9]), .C(R14[9]), .D(R15[9]), .S0(n988), 
        .S1(n996), .Y(n960) );
  MXI4X1 U1945 ( .A(R4[9]), .B(R5[9]), .C(R6[9]), .D(R7[9]), .S0(n988), .S1(
        n996), .Y(n959) );
  MXI4X1 U1946 ( .A(R8[9]), .B(R9[9]), .C(R10[9]), .D(R11[9]), .S0(n988), .S1(
        n996), .Y(n958) );
  MXI4X1 U1947 ( .A(n961), .B(n962), .C(n963), .D(n964), .S0(N56), .S1(N55), 
        .Y(N72) );
  MXI4X1 U1948 ( .A(R12[10]), .B(R13[10]), .C(R14[10]), .D(R15[10]), .S0(n989), 
        .S1(n997), .Y(n964) );
  MXI4X1 U1949 ( .A(R4[10]), .B(R5[10]), .C(R6[10]), .D(R7[10]), .S0(n989), 
        .S1(n997), .Y(n963) );
  MXI4X1 U1950 ( .A(R8[10]), .B(R9[10]), .C(R10[10]), .D(R11[10]), .S0(n989), 
        .S1(n997), .Y(n962) );
  MXI4X1 U1951 ( .A(n965), .B(n966), .C(n967), .D(n968), .S0(N56), .S1(N55), 
        .Y(N71) );
  MXI4X1 U1952 ( .A(R12[11]), .B(R13[11]), .C(R14[11]), .D(R15[11]), .S0(n989), 
        .S1(n997), .Y(n968) );
  MXI4X1 U1953 ( .A(R4[11]), .B(R5[11]), .C(R6[11]), .D(R7[11]), .S0(n989), 
        .S1(n997), .Y(n967) );
  MXI4X1 U1954 ( .A(R8[11]), .B(R9[11]), .C(R10[11]), .D(R11[11]), .S0(n989), 
        .S1(n997), .Y(n966) );
  MXI4X1 U1955 ( .A(n969), .B(n970), .C(n971), .D(n972), .S0(N56), .S1(N55), 
        .Y(N70) );
  MXI4X1 U1956 ( .A(R12[12]), .B(R13[12]), .C(R14[12]), .D(R15[12]), .S0(n989), 
        .S1(n997), .Y(n972) );
  MXI4X1 U1957 ( .A(R4[12]), .B(R5[12]), .C(R6[12]), .D(R7[12]), .S0(n989), 
        .S1(n997), .Y(n971) );
  MXI4X1 U1958 ( .A(R8[12]), .B(R9[12]), .C(R10[12]), .D(R11[12]), .S0(n989), 
        .S1(n997), .Y(n970) );
  MXI4X1 U1959 ( .A(n973), .B(n974), .C(n975), .D(n976), .S0(N56), .S1(N55), 
        .Y(N69) );
  MXI4X1 U1960 ( .A(R12[13]), .B(R13[13]), .C(R14[13]), .D(R15[13]), .S0(n990), 
        .S1(n998), .Y(n976) );
  MXI4X1 U1961 ( .A(R4[13]), .B(R5[13]), .C(R6[13]), .D(R7[13]), .S0(n990), 
        .S1(n998), .Y(n975) );
  MXI4X1 U1962 ( .A(R8[13]), .B(R9[13]), .C(R10[13]), .D(R11[13]), .S0(n990), 
        .S1(n998), .Y(n974) );
  MXI4X1 U1963 ( .A(n977), .B(n978), .C(n979), .D(n980), .S0(N56), .S1(N55), 
        .Y(N68) );
  MXI4X1 U1964 ( .A(R12[14]), .B(R13[14]), .C(R14[14]), .D(R15[14]), .S0(n990), 
        .S1(n998), .Y(n980) );
  MXI4X1 U1965 ( .A(R4[14]), .B(R5[14]), .C(R6[14]), .D(R7[14]), .S0(n990), 
        .S1(n998), .Y(n979) );
  MXI4X1 U1966 ( .A(R8[14]), .B(R9[14]), .C(R10[14]), .D(R11[14]), .S0(n990), 
        .S1(n998), .Y(n978) );
  MXI4X1 U1967 ( .A(n981), .B(n982), .C(n983), .D(n984), .S0(N56), .S1(N55), 
        .Y(N67) );
  MXI4X1 U1968 ( .A(R4[15]), .B(R5[15]), .C(R6[15]), .D(R7[15]), .S0(n990), 
        .S1(n998), .Y(n983) );
  MXI4X1 U1969 ( .A(R12[15]), .B(R13[15]), .C(R14[15]), .D(R15[15]), .S0(n990), 
        .S1(n998), .Y(n984) );
  MXI4X1 U1970 ( .A(R0[15]), .B(R1[15]), .C(R2[15]), .D(R3[15]), .S0(n990), 
        .S1(n998), .Y(n981) );
  MXI4X1 U1971 ( .A(R4[0]), .B(R5[0]), .C(R6[0]), .D(R7[0]), .S0(n985), .S1(
        n993), .Y(n923) );
  MXI4X1 U1972 ( .A(R4[1]), .B(R5[1]), .C(R6[1]), .D(R7[1]), .S0(n986), .S1(
        n994), .Y(n927) );
  MXI4X1 U1973 ( .A(R4[2]), .B(R5[2]), .C(R6[2]), .D(R7[2]), .S0(n986), .S1(
        n994), .Y(n931) );
  MXI4X1 U1974 ( .A(R4[3]), .B(R5[3]), .C(R6[3]), .D(R7[3]), .S0(n986), .S1(
        n994), .Y(n935) );
  MXI4X1 U1975 ( .A(R4[4]), .B(R5[4]), .C(R6[4]), .D(R7[4]), .S0(n987), .S1(
        n995), .Y(n939) );
  MXI4X1 U1976 ( .A(R4[5]), .B(R5[5]), .C(R6[5]), .D(R7[5]), .S0(n987), .S1(
        n995), .Y(n943) );
  MXI4X1 U1977 ( .A(R4[6]), .B(R5[6]), .C(R6[6]), .D(R7[6]), .S0(n987), .S1(
        n995), .Y(n947) );
  MXI4X1 U1978 ( .A(R4[7]), .B(R5[7]), .C(R6[7]), .D(R7[7]), .S0(n988), .S1(
        n996), .Y(n951) );
  MXI4X1 U1979 ( .A(R4[8]), .B(R5[8]), .C(R6[8]), .D(R7[8]), .S0(n988), .S1(
        n996), .Y(n955) );
  MXI4X1 U1980 ( .A(R0[0]), .B(R1[0]), .C(R2[0]), .D(R3[0]), .S0(n985), .S1(
        n993), .Y(n921) );
  MXI4X1 U1981 ( .A(R0[9]), .B(R1[9]), .C(R2[9]), .D(R3[9]), .S0(n988), .S1(
        n996), .Y(n957) );
  MXI4X1 U1982 ( .A(R0[10]), .B(R1[10]), .C(R2[10]), .D(R3[10]), .S0(n989), 
        .S1(n997), .Y(n961) );
  MXI4X1 U1983 ( .A(R0[11]), .B(R1[11]), .C(R2[11]), .D(R3[11]), .S0(n989), 
        .S1(n997), .Y(n965) );
  MXI4X1 U1984 ( .A(R0[12]), .B(R1[12]), .C(R2[12]), .D(R3[12]), .S0(n989), 
        .S1(n997), .Y(n969) );
  MXI4X1 U1985 ( .A(R0[13]), .B(R1[13]), .C(R2[13]), .D(R3[13]), .S0(n990), 
        .S1(n998), .Y(n973) );
  MXI4X1 U1986 ( .A(R0[14]), .B(R1[14]), .C(R2[14]), .D(R3[14]), .S0(n990), 
        .S1(n998), .Y(n977) );
  MXI4X1 U1987 ( .A(R0[1]), .B(R1[1]), .C(R2[1]), .D(R3[1]), .S0(n986), .S1(
        n994), .Y(n925) );
  MXI4X1 U1988 ( .A(R0[2]), .B(R1[2]), .C(R2[2]), .D(R3[2]), .S0(n986), .S1(
        n994), .Y(n929) );
  MXI4X1 U1989 ( .A(R0[3]), .B(R1[3]), .C(R2[3]), .D(R3[3]), .S0(n986), .S1(
        n994), .Y(n933) );
  MXI4X1 U1990 ( .A(R0[4]), .B(R1[4]), .C(R2[4]), .D(R3[4]), .S0(n987), .S1(
        n995), .Y(n937) );
  MXI4X1 U1991 ( .A(R0[5]), .B(R1[5]), .C(R2[5]), .D(R3[5]), .S0(n987), .S1(
        n995), .Y(n941) );
  MXI4X1 U1992 ( .A(R0[6]), .B(R1[6]), .C(R2[6]), .D(R3[6]), .S0(n987), .S1(
        n995), .Y(n945) );
  MXI4X1 U1993 ( .A(R0[7]), .B(R1[7]), .C(R2[7]), .D(R3[7]), .S0(n988), .S1(
        n996), .Y(n949) );
  MXI4X1 U1994 ( .A(R0[8]), .B(R1[8]), .C(R2[8]), .D(R3[8]), .S0(n988), .S1(
        n996), .Y(n953) );
  MXI4X1 U1995 ( .A(R8[0]), .B(R9[0]), .C(R10[0]), .D(R11[0]), .S0(n985), .S1(
        n993), .Y(n922) );
  MXI4X1 U1996 ( .A(R8[15]), .B(R9[15]), .C(R10[15]), .D(R11[15]), .S0(n990), 
        .S1(n998), .Y(n982) );
  MXI4X1 U1997 ( .A(R8[1]), .B(R9[1]), .C(R10[1]), .D(R11[1]), .S0(n986), .S1(
        n994), .Y(n926) );
  MXI4X1 U1998 ( .A(R8[2]), .B(R9[2]), .C(R10[2]), .D(R11[2]), .S0(n986), .S1(
        n994), .Y(n930) );
  MXI4X1 U1999 ( .A(R8[3]), .B(R9[3]), .C(R10[3]), .D(R11[3]), .S0(n986), .S1(
        n994), .Y(n934) );
  MXI4X1 U2000 ( .A(R8[4]), .B(R9[4]), .C(R10[4]), .D(R11[4]), .S0(n987), .S1(
        n995), .Y(n938) );
  MXI4X1 U2001 ( .A(R8[5]), .B(R9[5]), .C(R10[5]), .D(R11[5]), .S0(n987), .S1(
        n995), .Y(n942) );
  MXI4X1 U2002 ( .A(R8[6]), .B(R9[6]), .C(R10[6]), .D(R11[6]), .S0(n987), .S1(
        n995), .Y(n946) );
  MXI4X1 U2003 ( .A(R8[7]), .B(R9[7]), .C(R10[7]), .D(R11[7]), .S0(n988), .S1(
        n996), .Y(n950) );
  MXI4X1 U2004 ( .A(R8[8]), .B(R9[8]), .C(R10[8]), .D(R11[8]), .S0(n988), .S1(
        n996), .Y(n954) );
  NOR2BX1 U2005 ( .AN(control[1]), .B(n1868), .Y(n129) );
  NOR2X1 U2006 ( .A(n1868), .B(control[1]), .Y(n128) );
  NOR2X1 U2007 ( .A(n1831), .B(n1714), .Y(n1715) );
  CLKINVX1 U2008 ( .A(data[9]), .Y(n1714) );
  NOR2X1 U2009 ( .A(n1831), .B(n1750), .Y(n1751) );
  CLKINVX1 U2010 ( .A(data[11]), .Y(n1750) );
  NOR2X1 U2011 ( .A(n1831), .B(n1787), .Y(n1788) );
  CLKINVX1 U2012 ( .A(data[13]), .Y(n1787) );
  CLKINVX1 U2013 ( .A(N55), .Y(n1867) );
  CLKINVX1 U2014 ( .A(N56), .Y(n1866) );
  CLKBUFX3 U2015 ( .A(N54), .Y(n1000) );
  CLKBUFX3 U2016 ( .A(N54), .Y(n999) );
  CLKINVX1 U2017 ( .A(data[10]), .Y(n1732) );
  CLKINVX1 U2018 ( .A(data[12]), .Y(n1770) );
  CLKINVX1 U2019 ( .A(data[14]), .Y(n1808) );
  CLKINVX1 U2020 ( .A(data[15]), .Y(n1830) );
  NAND3X1 U2021 ( .A(n1744), .B(n1743), .C(n1742), .Y(n1780) );
  NAND2X1 U2022 ( .A(n1173), .B(n1744), .Y(n1721) );
  NAND2X1 U2023 ( .A(\add_233/carry[6] ), .B(n1173), .Y(n1656) );
  AOI2BB2X2 U2024 ( .B0(N528), .B1(n1852), .A0N(n1811), .A1N(n1810), .Y(n1829)
         );
  OAI21XL U2025 ( .A0(\add_233/carry[8] ), .A1(n1814), .B0(n1687), .Y(n1692)
         );
  NOR2X1 U2026 ( .A(n1864), .B(n1863), .Y(V) );
  OR2X1 U2027 ( .A(BUSA[6]), .B(\add_233/carry[6] ), .Y(\add_233/carry[7] ) );
  OR2X1 U2028 ( .A(BUSA[3]), .B(\add_233/carry[3] ), .Y(\add_233/carry[4] ) );
  OR2X1 U2029 ( .A(BUSA[2]), .B(\add_233/carry[2] ), .Y(\add_233/carry[3] ) );
endmodule

